-- DUAL_PORT_RAM.vhd