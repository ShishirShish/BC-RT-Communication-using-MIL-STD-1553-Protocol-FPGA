`timescale 1 ns/100 ps
// Version: 2025.2 2025.2.0.14


module bcrt(
       FIC_0_ACLK,
       FIC_0_AXI4_M_AWREADY,
       FIC_0_AXI4_M_WREADY,
       FIC_0_AXI4_M_BID,
       FIC_0_AXI4_M_BRESP,
       FIC_0_AXI4_M_BVALID,
       FIC_0_AXI4_M_ARREADY,
       FIC_0_AXI4_M_RID,
       FIC_0_AXI4_M_RDATA,
       FIC_0_AXI4_M_RRESP,
       FIC_0_AXI4_M_RLAST,
       FIC_0_AXI4_M_RVALID,
       FIC_0_AXI4_S_AWID,
       FIC_0_AXI4_S_AWADDR,
       FIC_0_AXI4_S_AWLEN,
       FIC_0_AXI4_S_AWSIZE,
       FIC_0_AXI4_S_AWBURST,
       FIC_0_AXI4_S_AWQOS,
       FIC_0_AXI4_S_AWLOCK,
       FIC_0_AXI4_S_AWCACHE,
       FIC_0_AXI4_S_AWPROT,
       FIC_0_AXI4_S_AWVALID,
       FIC_0_AXI4_S_WDATA,
       FIC_0_AXI4_S_WSTRB,
       FIC_0_AXI4_S_WLAST,
       FIC_0_AXI4_S_WVALID,
       FIC_0_AXI4_S_BREADY,
       FIC_0_AXI4_S_ARID,
       FIC_0_AXI4_S_ARADDR,
       FIC_0_AXI4_S_ARLEN,
       FIC_0_AXI4_S_ARSIZE,
       FIC_0_AXI4_S_ARBURST,
       FIC_0_AXI4_S_ARQOS,
       FIC_0_AXI4_S_ARLOCK,
       FIC_0_AXI4_S_ARCACHE,
       FIC_0_AXI4_S_ARPROT,
       FIC_0_AXI4_S_ARVALID,
       FIC_0_AXI4_S_RREADY,
       FIC_1_ACLK,
       FIC_1_AXI4_S_AWID,
       FIC_1_AXI4_S_AWADDR,
       FIC_1_AXI4_S_AWLEN,
       FIC_1_AXI4_S_AWSIZE,
       FIC_1_AXI4_S_AWBURST,
       FIC_1_AXI4_S_AWLOCK,
       FIC_1_AXI4_S_AWCACHE,
       FIC_1_AXI4_S_AWQOS,
       FIC_1_AXI4_S_AWPROT,
       FIC_1_AXI4_S_AWVALID,
       FIC_1_AXI4_S_WDATA,
       FIC_1_AXI4_S_WSTRB,
       FIC_1_AXI4_S_WLAST,
       FIC_1_AXI4_S_WVALID,
       FIC_1_AXI4_S_BREADY,
       FIC_1_AXI4_S_ARID,
       FIC_1_AXI4_S_ARADDR,
       FIC_1_AXI4_S_ARLEN,
       FIC_1_AXI4_S_ARSIZE,
       FIC_1_AXI4_S_ARBURST,
       FIC_1_AXI4_S_ARQOS,
       FIC_1_AXI4_S_ARLOCK,
       FIC_1_AXI4_S_ARCACHE,
       FIC_1_AXI4_S_ARPROT,
       FIC_1_AXI4_S_ARVALID,
       FIC_1_AXI4_S_RREADY,
       FIC_2_ACLK,
       FIC_2_AXI4_S_AWID,
       FIC_2_AXI4_S_AWADDR,
       FIC_2_AXI4_S_AWLEN,
       FIC_2_AXI4_S_AWSIZE,
       FIC_2_AXI4_S_AWBURST,
       FIC_2_AXI4_S_AWLOCK,
       FIC_2_AXI4_S_AWCACHE,
       FIC_2_AXI4_S_AWQOS,
       FIC_2_AXI4_S_AWPROT,
       FIC_2_AXI4_S_AWVALID,
       FIC_2_AXI4_S_WDATA,
       FIC_2_AXI4_S_WSTRB,
       FIC_2_AXI4_S_WLAST,
       FIC_2_AXI4_S_WVALID,
       FIC_2_AXI4_S_BREADY,
       FIC_2_AXI4_S_ARID,
       FIC_2_AXI4_S_ARADDR,
       FIC_2_AXI4_S_ARLEN,
       FIC_2_AXI4_S_ARSIZE,
       FIC_2_AXI4_S_ARBURST,
       FIC_2_AXI4_S_ARLOCK,
       FIC_2_AXI4_S_ARCACHE,
       FIC_2_AXI4_S_ARQOS,
       FIC_2_AXI4_S_ARPROT,
       FIC_2_AXI4_S_ARVALID,
       FIC_2_AXI4_S_RREADY,
       FIC_3_PCLK,
       FIC_3_APB_M_PRDATA,
       FIC_3_APB_M_PREADY,
       FIC_3_APB_M_PSLVERR,
       MMUART_0_RXD_F2M,
       MMUART_1_RXD_F2M,
       MMUART_2_RXD_F2M,
       MMUART_3_RXD_F2M,
       MMUART_4_RXD_F2M,
       CAN_0_RXBUS_F2M,
       QSPI_DATA2_F2M,
       QSPI_DATA3_F2M,
       SPI_0_SS_F2M,
       SPI_0_DI_F2M,
       SPI_0_CLK_F2M,
       I2C_0_SCL_F2M,
       I2C_0_SDA_F2M,
       GPIO_2_F2M_31,
       GPIO_2_F2M_30,
       MSS_INT_F2M,
       MSS_RESET_N_F2M,
       FIC_0_DLL_LOCK_M2F,
       FIC_1_DLL_LOCK_M2F,
       FIC_2_DLL_LOCK_M2F,
       FIC_3_DLL_LOCK_M2F,
       FIC_0_AXI4_M_AWID,
       FIC_0_AXI4_M_AWADDR,
       FIC_0_AXI4_M_AWLEN,
       FIC_0_AXI4_M_AWSIZE,
       FIC_0_AXI4_M_AWBURST,
       FIC_0_AXI4_M_AWLOCK,
       FIC_0_AXI4_M_AWQOS,
       FIC_0_AXI4_M_AWCACHE,
       FIC_0_AXI4_M_AWPROT,
       FIC_0_AXI4_M_AWVALID,
       FIC_0_AXI4_M_WDATA,
       FIC_0_AXI4_M_WSTRB,
       FIC_0_AXI4_M_WLAST,
       FIC_0_AXI4_M_WVALID,
       FIC_0_AXI4_M_BREADY,
       FIC_0_AXI4_M_ARID,
       FIC_0_AXI4_M_ARADDR,
       FIC_0_AXI4_M_ARLEN,
       FIC_0_AXI4_M_ARSIZE,
       FIC_0_AXI4_M_ARBURST,
       FIC_0_AXI4_M_ARLOCK,
       FIC_0_AXI4_M_ARQOS,
       FIC_0_AXI4_M_ARCACHE,
       FIC_0_AXI4_M_ARPROT,
       FIC_0_AXI4_M_ARVALID,
       FIC_0_AXI4_M_RREADY,
       FIC_0_AXI4_S_AWREADY,
       FIC_0_AXI4_S_WREADY,
       FIC_0_AXI4_S_BID,
       FIC_0_AXI4_S_BRESP,
       FIC_0_AXI4_S_BVALID,
       FIC_0_AXI4_S_ARREADY,
       FIC_0_AXI4_S_RID,
       FIC_0_AXI4_S_RDATA,
       FIC_0_AXI4_S_RRESP,
       FIC_0_AXI4_S_RLAST,
       FIC_0_AXI4_S_RVALID,
       FIC_1_AXI4_S_AWREADY,
       FIC_1_AXI4_S_WREADY,
       FIC_1_AXI4_S_BID,
       FIC_1_AXI4_S_BRESP,
       FIC_1_AXI4_S_BVALID,
       FIC_1_AXI4_S_ARREADY,
       FIC_1_AXI4_S_RID,
       FIC_1_AXI4_S_RDATA,
       FIC_1_AXI4_S_RRESP,
       FIC_1_AXI4_S_RLAST,
       FIC_1_AXI4_S_RVALID,
       FIC_2_AXI4_S_AWREADY,
       FIC_2_AXI4_S_WREADY,
       FIC_2_AXI4_S_BID,
       FIC_2_AXI4_S_BRESP,
       FIC_2_AXI4_S_BVALID,
       FIC_2_AXI4_S_ARREADY,
       FIC_2_AXI4_S_RID,
       FIC_2_AXI4_S_RDATA,
       FIC_2_AXI4_S_RRESP,
       FIC_2_AXI4_S_RLAST,
       FIC_2_AXI4_S_RVALID,
       FIC_3_APB_M_PSEL,
       FIC_3_APB_M_PADDR,
       FIC_3_APB_M_PWRITE,
       FIC_3_APB_M_PENABLE,
       FIC_3_APB_M_PSTRB,
       FIC_3_APB_M_PWDATA,
       MMUART_0_TXD_M2F,
       MMUART_0_TXD_OE_M2F,
       MMUART_1_TXD_M2F,
       MMUART_1_TXD_OE_M2F,
       MMUART_2_TXD_M2F,
       MMUART_3_TXD_M2F,
       MMUART_4_TXD_M2F,
       CAN_0_TX_EBL_M2F,
       CAN_0_TXBUS_M2F,
       QSPI_DATA2_M2F,
       QSPI_DATA3_M2F,
       QSPI_DATA2_OE_M2F,
       QSPI_DATA3_OE_M2F,
       SPI_0_SS1_M2F,
       SPI_0_SS1_OE_M2F,
       SPI_0_DO_M2F,
       SPI_0_DO_OE_M2F,
       SPI_0_CLK_M2F,
       SPI_0_CLK_OE_M2F,
       I2C_0_SCL_OE_M2F,
       I2C_0_SDA_OE_M2F,
       GPIO_2_M2F_28,
       GPIO_2_M2F_27,
       GPIO_2_M2F_26,
       GPIO_2_M2F_19,
       GPIO_2_M2F_18,
       GPIO_2_M2F_17,
       GPIO_2_M2F_16,
       MSS_INT_M2F,
       PLL_CPU_LOCK_M2F,
       PLL_DDR_LOCK_M2F,
       PLL_SGMII_LOCK_M2F,
       MSS_RESET_N_M2F,
       MAC_0_TSU_SOF_TX_M2F,
       MAC_0_TSU_SYNC_FRAME_TX_M2F,
       MAC_0_TSU_DELAY_REQ_TX_M2F,
       MAC_0_TSU_PDELAY_REQ_TX_M2F,
       MAC_0_TSU_PDELAY_RESP_TX_M2F,
       MAC_0_TSU_SOF_RX_M2F,
       MAC_0_TSU_SYNC_FRAME_RX_M2F,
       MAC_0_TSU_DELAY_REQ_RX_M2F,
       MAC_0_TSU_PDELAY_REQ_RX_M2F,
       MAC_0_TSU_PDELAY_RESP_RX_M2F,
       MAC_0_TSU_TIMER_CNT_M2F,
       MAC_1_TSU_SOF_TX_M2F,
       MAC_1_TSU_SYNC_FRAME_TX_M2F,
       MAC_1_TSU_DELAY_REQ_TX_M2F,
       MAC_1_TSU_PDELAY_REQ_TX_M2F,
       MAC_1_TSU_PDELAY_RESP_TX_M2F,
       MAC_1_TSU_SOF_RX_M2F,
       MAC_1_TSU_SYNC_FRAME_RX_M2F,
       MAC_1_TSU_DELAY_REQ_RX_M2F,
       MAC_1_TSU_PDELAY_REQ_RX_M2F,
       MAC_1_TSU_PDELAY_RESP_RX_M2F,
       MAC_1_TSU_TIMER_CNT_M2F,
       I2C_1_SCL,
       I2C_1_SDA,
       CAN_1_TXBUS,
       CAN_1_RXBUS,
       CAN_1_TX_EBL_N,
       MAC_1_MDIO,
       MAC_1_MDC,
       USB_CLK,
       USB_DIR,
       USB_NXT,
       USB_STP,
       USB_DATA0,
       USB_DATA1,
       USB_DATA2,
       USB_DATA3,
       USB_DATA4,
       USB_DATA5,
       USB_DATA6,
       USB_DATA7,
       QSPI_DATA0,
       QSPI_DATA1,
       QSPI_SS0,
       QSPI_CLK,
       EMMC_CLK_SD_CLK,
       EMMC_CMD_SD_CMD,
       EMMC_DATA0_SD_DATA0,
       EMMC_DATA1_SD_DATA1,
       EMMC_DATA2_SD_DATA2,
       EMMC_DATA3_SD_DATA3,
       EMMC_DATA4_SD_POW,
       EMMC_DATA5_SD_VOLT_SEL,
       EMMC_DATA6_SD_VOLT_EN,
       EMMC_DATA7_SD_VOLT_CMD_DIR,
       EMMC_UNUSED_SD_VOLT_DIR_0,
       EMMC_UNUSED_SD_VOLT_DIR_1_3,
       EMMC_STRB_SD_CD,
       EMMC_RSTN_SD_WP,
       SGMII_RX1_P,
       SGMII_RX1_N,
       SGMII_RX0_P,
       SGMII_RX0_N,
       SGMII_TX1_P,
       SGMII_TX1_N,
       SGMII_TX0_P,
       SGMII_TX0_N,
       REFCLK,
       REFCLK_N,
       DQ,
       DQS,
       DQS_N,
       DM,
       RESET_N,
       ODT,
       CKE,
       CS,
       CK,
       CK_N,
       CA
    );
input  FIC_0_ACLK;
input  FIC_0_AXI4_M_AWREADY;
input  FIC_0_AXI4_M_WREADY;
input  [7:0] FIC_0_AXI4_M_BID;
input  [1:0] FIC_0_AXI4_M_BRESP;
input  FIC_0_AXI4_M_BVALID;
input  FIC_0_AXI4_M_ARREADY;
input  [7:0] FIC_0_AXI4_M_RID;
input  [63:0] FIC_0_AXI4_M_RDATA;
input  [1:0] FIC_0_AXI4_M_RRESP;
input  FIC_0_AXI4_M_RLAST;
input  FIC_0_AXI4_M_RVALID;
input  [3:0] FIC_0_AXI4_S_AWID;
input  [37:0] FIC_0_AXI4_S_AWADDR;
input  [7:0] FIC_0_AXI4_S_AWLEN;
input  [2:0] FIC_0_AXI4_S_AWSIZE;
input  [1:0] FIC_0_AXI4_S_AWBURST;
input  [3:0] FIC_0_AXI4_S_AWQOS;
input  FIC_0_AXI4_S_AWLOCK;
input  [3:0] FIC_0_AXI4_S_AWCACHE;
input  [2:0] FIC_0_AXI4_S_AWPROT;
input  FIC_0_AXI4_S_AWVALID;
input  [63:0] FIC_0_AXI4_S_WDATA;
input  [7:0] FIC_0_AXI4_S_WSTRB;
input  FIC_0_AXI4_S_WLAST;
input  FIC_0_AXI4_S_WVALID;
input  FIC_0_AXI4_S_BREADY;
input  [3:0] FIC_0_AXI4_S_ARID;
input  [37:0] FIC_0_AXI4_S_ARADDR;
input  [7:0] FIC_0_AXI4_S_ARLEN;
input  [2:0] FIC_0_AXI4_S_ARSIZE;
input  [1:0] FIC_0_AXI4_S_ARBURST;
input  [3:0] FIC_0_AXI4_S_ARQOS;
input  FIC_0_AXI4_S_ARLOCK;
input  [3:0] FIC_0_AXI4_S_ARCACHE;
input  [2:0] FIC_0_AXI4_S_ARPROT;
input  FIC_0_AXI4_S_ARVALID;
input  FIC_0_AXI4_S_RREADY;
input  FIC_1_ACLK;
input  [3:0] FIC_1_AXI4_S_AWID;
input  [37:0] FIC_1_AXI4_S_AWADDR;
input  [7:0] FIC_1_AXI4_S_AWLEN;
input  [2:0] FIC_1_AXI4_S_AWSIZE;
input  [1:0] FIC_1_AXI4_S_AWBURST;
input  FIC_1_AXI4_S_AWLOCK;
input  [3:0] FIC_1_AXI4_S_AWCACHE;
input  [3:0] FIC_1_AXI4_S_AWQOS;
input  [2:0] FIC_1_AXI4_S_AWPROT;
input  FIC_1_AXI4_S_AWVALID;
input  [63:0] FIC_1_AXI4_S_WDATA;
input  [7:0] FIC_1_AXI4_S_WSTRB;
input  FIC_1_AXI4_S_WLAST;
input  FIC_1_AXI4_S_WVALID;
input  FIC_1_AXI4_S_BREADY;
input  [3:0] FIC_1_AXI4_S_ARID;
input  [37:0] FIC_1_AXI4_S_ARADDR;
input  [7:0] FIC_1_AXI4_S_ARLEN;
input  [2:0] FIC_1_AXI4_S_ARSIZE;
input  [1:0] FIC_1_AXI4_S_ARBURST;
input  [3:0] FIC_1_AXI4_S_ARQOS;
input  FIC_1_AXI4_S_ARLOCK;
input  [3:0] FIC_1_AXI4_S_ARCACHE;
input  [2:0] FIC_1_AXI4_S_ARPROT;
input  FIC_1_AXI4_S_ARVALID;
input  FIC_1_AXI4_S_RREADY;
input  FIC_2_ACLK;
input  [3:0] FIC_2_AXI4_S_AWID;
input  [37:0] FIC_2_AXI4_S_AWADDR;
input  [7:0] FIC_2_AXI4_S_AWLEN;
input  [2:0] FIC_2_AXI4_S_AWSIZE;
input  [1:0] FIC_2_AXI4_S_AWBURST;
input  FIC_2_AXI4_S_AWLOCK;
input  [3:0] FIC_2_AXI4_S_AWCACHE;
input  [3:0] FIC_2_AXI4_S_AWQOS;
input  [2:0] FIC_2_AXI4_S_AWPROT;
input  FIC_2_AXI4_S_AWVALID;
input  [63:0] FIC_2_AXI4_S_WDATA;
input  [7:0] FIC_2_AXI4_S_WSTRB;
input  FIC_2_AXI4_S_WLAST;
input  FIC_2_AXI4_S_WVALID;
input  FIC_2_AXI4_S_BREADY;
input  [3:0] FIC_2_AXI4_S_ARID;
input  [37:0] FIC_2_AXI4_S_ARADDR;
input  [7:0] FIC_2_AXI4_S_ARLEN;
input  [2:0] FIC_2_AXI4_S_ARSIZE;
input  [1:0] FIC_2_AXI4_S_ARBURST;
input  FIC_2_AXI4_S_ARLOCK;
input  [3:0] FIC_2_AXI4_S_ARCACHE;
input  [3:0] FIC_2_AXI4_S_ARQOS;
input  [2:0] FIC_2_AXI4_S_ARPROT;
input  FIC_2_AXI4_S_ARVALID;
input  FIC_2_AXI4_S_RREADY;
input  FIC_3_PCLK;
input  [31:0] FIC_3_APB_M_PRDATA;
input  FIC_3_APB_M_PREADY;
input  FIC_3_APB_M_PSLVERR;
input  MMUART_0_RXD_F2M;
input  MMUART_1_RXD_F2M;
input  MMUART_2_RXD_F2M;
input  MMUART_3_RXD_F2M;
input  MMUART_4_RXD_F2M;
input  CAN_0_RXBUS_F2M;
input  QSPI_DATA2_F2M;
input  QSPI_DATA3_F2M;
input  SPI_0_SS_F2M;
input  SPI_0_DI_F2M;
input  SPI_0_CLK_F2M;
input  I2C_0_SCL_F2M;
input  I2C_0_SDA_F2M;
input  GPIO_2_F2M_31;
input  GPIO_2_F2M_30;
input  [63:0] MSS_INT_F2M;
input  MSS_RESET_N_F2M;
output FIC_0_DLL_LOCK_M2F;
output FIC_1_DLL_LOCK_M2F;
output FIC_2_DLL_LOCK_M2F;
output FIC_3_DLL_LOCK_M2F;
output [7:0] FIC_0_AXI4_M_AWID;
output [37:0] FIC_0_AXI4_M_AWADDR;
output [7:0] FIC_0_AXI4_M_AWLEN;
output [2:0] FIC_0_AXI4_M_AWSIZE;
output [1:0] FIC_0_AXI4_M_AWBURST;
output FIC_0_AXI4_M_AWLOCK;
output [3:0] FIC_0_AXI4_M_AWQOS;
output [3:0] FIC_0_AXI4_M_AWCACHE;
output [2:0] FIC_0_AXI4_M_AWPROT;
output FIC_0_AXI4_M_AWVALID;
output [63:0] FIC_0_AXI4_M_WDATA;
output [7:0] FIC_0_AXI4_M_WSTRB;
output FIC_0_AXI4_M_WLAST;
output FIC_0_AXI4_M_WVALID;
output FIC_0_AXI4_M_BREADY;
output [7:0] FIC_0_AXI4_M_ARID;
output [37:0] FIC_0_AXI4_M_ARADDR;
output [7:0] FIC_0_AXI4_M_ARLEN;
output [2:0] FIC_0_AXI4_M_ARSIZE;
output [1:0] FIC_0_AXI4_M_ARBURST;
output FIC_0_AXI4_M_ARLOCK;
output [3:0] FIC_0_AXI4_M_ARQOS;
output [3:0] FIC_0_AXI4_M_ARCACHE;
output [2:0] FIC_0_AXI4_M_ARPROT;
output FIC_0_AXI4_M_ARVALID;
output FIC_0_AXI4_M_RREADY;
output FIC_0_AXI4_S_AWREADY;
output FIC_0_AXI4_S_WREADY;
output [3:0] FIC_0_AXI4_S_BID;
output [1:0] FIC_0_AXI4_S_BRESP;
output FIC_0_AXI4_S_BVALID;
output FIC_0_AXI4_S_ARREADY;
output [3:0] FIC_0_AXI4_S_RID;
output [63:0] FIC_0_AXI4_S_RDATA;
output [1:0] FIC_0_AXI4_S_RRESP;
output FIC_0_AXI4_S_RLAST;
output FIC_0_AXI4_S_RVALID;
output FIC_1_AXI4_S_AWREADY;
output FIC_1_AXI4_S_WREADY;
output [3:0] FIC_1_AXI4_S_BID;
output [1:0] FIC_1_AXI4_S_BRESP;
output FIC_1_AXI4_S_BVALID;
output FIC_1_AXI4_S_ARREADY;
output [3:0] FIC_1_AXI4_S_RID;
output [63:0] FIC_1_AXI4_S_RDATA;
output [1:0] FIC_1_AXI4_S_RRESP;
output FIC_1_AXI4_S_RLAST;
output FIC_1_AXI4_S_RVALID;
output FIC_2_AXI4_S_AWREADY;
output FIC_2_AXI4_S_WREADY;
output [3:0] FIC_2_AXI4_S_BID;
output [1:0] FIC_2_AXI4_S_BRESP;
output FIC_2_AXI4_S_BVALID;
output FIC_2_AXI4_S_ARREADY;
output [3:0] FIC_2_AXI4_S_RID;
output [63:0] FIC_2_AXI4_S_RDATA;
output [1:0] FIC_2_AXI4_S_RRESP;
output FIC_2_AXI4_S_RLAST;
output FIC_2_AXI4_S_RVALID;
output FIC_3_APB_M_PSEL;
output [31:0] FIC_3_APB_M_PADDR;
output FIC_3_APB_M_PWRITE;
output FIC_3_APB_M_PENABLE;
output [3:0] FIC_3_APB_M_PSTRB;
output [31:0] FIC_3_APB_M_PWDATA;
output MMUART_0_TXD_M2F;
output MMUART_0_TXD_OE_M2F;
output MMUART_1_TXD_M2F;
output MMUART_1_TXD_OE_M2F;
output MMUART_2_TXD_M2F;
output MMUART_3_TXD_M2F;
output MMUART_4_TXD_M2F;
output CAN_0_TX_EBL_M2F;
output CAN_0_TXBUS_M2F;
output QSPI_DATA2_M2F;
output QSPI_DATA3_M2F;
output QSPI_DATA2_OE_M2F;
output QSPI_DATA3_OE_M2F;
output SPI_0_SS1_M2F;
output SPI_0_SS1_OE_M2F;
output SPI_0_DO_M2F;
output SPI_0_DO_OE_M2F;
output SPI_0_CLK_M2F;
output SPI_0_CLK_OE_M2F;
output I2C_0_SCL_OE_M2F;
output I2C_0_SDA_OE_M2F;
output GPIO_2_M2F_28;
output GPIO_2_M2F_27;
output GPIO_2_M2F_26;
output GPIO_2_M2F_19;
output GPIO_2_M2F_18;
output GPIO_2_M2F_17;
output GPIO_2_M2F_16;
output [15:0] MSS_INT_M2F;
output PLL_CPU_LOCK_M2F;
output PLL_DDR_LOCK_M2F;
output PLL_SGMII_LOCK_M2F;
output MSS_RESET_N_M2F;
output MAC_0_TSU_SOF_TX_M2F;
output MAC_0_TSU_SYNC_FRAME_TX_M2F;
output MAC_0_TSU_DELAY_REQ_TX_M2F;
output MAC_0_TSU_PDELAY_REQ_TX_M2F;
output MAC_0_TSU_PDELAY_RESP_TX_M2F;
output MAC_0_TSU_SOF_RX_M2F;
output MAC_0_TSU_SYNC_FRAME_RX_M2F;
output MAC_0_TSU_DELAY_REQ_RX_M2F;
output MAC_0_TSU_PDELAY_REQ_RX_M2F;
output MAC_0_TSU_PDELAY_RESP_RX_M2F;
output [93:0] MAC_0_TSU_TIMER_CNT_M2F;
output MAC_1_TSU_SOF_TX_M2F;
output MAC_1_TSU_SYNC_FRAME_TX_M2F;
output MAC_1_TSU_DELAY_REQ_TX_M2F;
output MAC_1_TSU_PDELAY_REQ_TX_M2F;
output MAC_1_TSU_PDELAY_RESP_TX_M2F;
output MAC_1_TSU_SOF_RX_M2F;
output MAC_1_TSU_SYNC_FRAME_RX_M2F;
output MAC_1_TSU_DELAY_REQ_RX_M2F;
output MAC_1_TSU_PDELAY_REQ_RX_M2F;
output MAC_1_TSU_PDELAY_RESP_RX_M2F;
output [93:0] MAC_1_TSU_TIMER_CNT_M2F;
inout  I2C_1_SCL;
inout  I2C_1_SDA;
output CAN_1_TXBUS;
input  CAN_1_RXBUS;
output CAN_1_TX_EBL_N;
inout  MAC_1_MDIO;
output MAC_1_MDC;
input  USB_CLK;
input  USB_DIR;
input  USB_NXT;
output USB_STP;
inout  USB_DATA0;
inout  USB_DATA1;
inout  USB_DATA2;
inout  USB_DATA3;
inout  USB_DATA4;
inout  USB_DATA5;
inout  USB_DATA6;
inout  USB_DATA7;
inout  QSPI_DATA0;
inout  QSPI_DATA1;
output QSPI_SS0;
output QSPI_CLK;
output EMMC_CLK_SD_CLK;
inout  EMMC_CMD_SD_CMD;
inout  EMMC_DATA0_SD_DATA0;
inout  EMMC_DATA1_SD_DATA1;
inout  EMMC_DATA2_SD_DATA2;
inout  EMMC_DATA3_SD_DATA3;
inout  EMMC_DATA4_SD_POW;
inout  EMMC_DATA5_SD_VOLT_SEL;
inout  EMMC_DATA6_SD_VOLT_EN;
inout  EMMC_DATA7_SD_VOLT_CMD_DIR;
output EMMC_UNUSED_SD_VOLT_DIR_0;
output EMMC_UNUSED_SD_VOLT_DIR_1_3;
input  EMMC_STRB_SD_CD;
output EMMC_RSTN_SD_WP;
input  SGMII_RX1_P;
input  SGMII_RX1_N;
input  SGMII_RX0_P;
input  SGMII_RX0_N;
output SGMII_TX1_P;
output SGMII_TX1_N;
output SGMII_TX0_P;
output SGMII_TX0_N;
input  REFCLK;
input  REFCLK_N;
inout  [15:0] DQ;
inout  [1:0] DQS;
inout  [1:0] DQS_N;
output [1:0] DM;
output RESET_N;
output ODT;
output CKE;
output CS;
output CK;
output CK_N;
output [5:0] CA;

    wire GND_net, I2C_0_SCL_OE_M2F_I_MSS_net, 
        I2C_0_SDA_OE_M2F_I_MSS_net, D_MSSIO26_OUT_IOINST_net, 
        E_MSSIO26_OUT_IOINST_net, Y_MSSIO26_OUT_IOINST_net, 
        D_MSSIO27_OUT_IOINST_net, E_MSSIO27_OUT_IOINST_net, 
        Y_MSSIO27_OUT_IOINST_net, D_MSSIO34_OUT_IOINST_net, 
        Y_MSSIO35_IN_IOINST_net, D_MSSIO36_OUT_IOINST_net, 
        D_MSSIO29_OUT_IOINST_net, E_MSSIO29_OUT_IOINST_net, 
        Y_MSSIO29_OUT_IOINST_net, D_MSSIO28_OUT_IOINST_net, 
        Y_MSSIO14_IN_IOINST_net, Y_MSSIO15_IN_IOINST_net, 
        Y_MSSIO16_IN_IOINST_net, D_MSSIO17_OUT_IOINST_net, 
        D_MSSIO18_OUT_IOINST_net, E_MSSIO18_OUT_IOINST_net, 
        Y_MSSIO18_OUT_IOINST_net, D_MSSIO19_OUT_IOINST_net, 
        E_MSSIO19_OUT_IOINST_net, Y_MSSIO19_OUT_IOINST_net, 
        D_MSSIO20_OUT_IOINST_net, E_MSSIO20_OUT_IOINST_net, 
        Y_MSSIO20_OUT_IOINST_net, D_MSSIO21_OUT_IOINST_net, 
        E_MSSIO21_OUT_IOINST_net, Y_MSSIO21_OUT_IOINST_net, 
        D_MSSIO22_OUT_IOINST_net, E_MSSIO22_OUT_IOINST_net, 
        Y_MSSIO22_OUT_IOINST_net, D_MSSIO23_OUT_IOINST_net, 
        E_MSSIO23_OUT_IOINST_net, Y_MSSIO23_OUT_IOINST_net, 
        D_MSSIO24_OUT_IOINST_net, E_MSSIO24_OUT_IOINST_net, 
        Y_MSSIO24_OUT_IOINST_net, D_MSSIO25_OUT_IOINST_net, 
        E_MSSIO25_OUT_IOINST_net, Y_MSSIO25_OUT_IOINST_net, 
        D_MSSIO32_OUT_IOINST_net, E_MSSIO32_OUT_IOINST_net, 
        Y_MSSIO32_OUT_IOINST_net, D_MSSIO33_OUT_IOINST_net, 
        E_MSSIO33_OUT_IOINST_net, Y_MSSIO33_OUT_IOINST_net, 
        D_MSSIO31_OUT_IOINST_net, D_MSSIO30_OUT_IOINST_net, 
        D_MSSIO0_OUT_IOINST_net, D_MSSIO1_OUT_IOINST_net, 
        E_MSSIO1_OUT_IOINST_net, Y_MSSIO1_OUT_IOINST_net, 
        D_MSSIO2_OUT_IOINST_net, E_MSSIO2_OUT_IOINST_net, 
        Y_MSSIO2_OUT_IOINST_net, D_MSSIO3_OUT_IOINST_net, 
        E_MSSIO3_OUT_IOINST_net, Y_MSSIO3_OUT_IOINST_net, 
        D_MSSIO4_OUT_IOINST_net, E_MSSIO4_OUT_IOINST_net, 
        Y_MSSIO4_OUT_IOINST_net, D_MSSIO5_OUT_IOINST_net, 
        E_MSSIO5_OUT_IOINST_net, Y_MSSIO5_OUT_IOINST_net, 
        D_MSSIO8_OUT_IOINST_net, E_MSSIO8_OUT_IOINST_net, 
        Y_MSSIO8_OUT_IOINST_net, D_MSSIO9_OUT_IOINST_net, 
        E_MSSIO9_OUT_IOINST_net, Y_MSSIO9_OUT_IOINST_net, 
        D_MSSIO10_OUT_IOINST_net, E_MSSIO10_OUT_IOINST_net, 
        Y_MSSIO10_OUT_IOINST_net, D_MSSIO11_OUT_IOINST_net, 
        E_MSSIO11_OUT_IOINST_net, Y_MSSIO11_OUT_IOINST_net, 
        D_MSSIO12_OUT_IOINST_net, D_MSSIO13_OUT_IOINST_net, 
        Y_MSSIO6_IN_IOINST_net, D_MSSIO7_OUT_IOINST_net, 
        Y_SGMII_RX1_IOINST_net, Y_SGMII_RX0_IOINST_net, 
        D_SGMII_TX1_IOINST_net, D_SGMII_TX0_IOINST_net, 
        Y_REFCLK_IOINST_net, D_DDR_DQ15_OUT_IOINST_net, 
        E_DDR_DQ15_OUT_IOINST_net, Y_DDR_DQ15_OUT_IOINST_net, 
        D_DDR_DQ14_OUT_IOINST_net, E_DDR_DQ14_OUT_IOINST_net, 
        Y_DDR_DQ14_OUT_IOINST_net, D_DDR_DQ13_OUT_IOINST_net, 
        E_DDR_DQ13_OUT_IOINST_net, Y_DDR_DQ13_OUT_IOINST_net, 
        D_DDR_DQ12_OUT_IOINST_net, E_DDR_DQ12_OUT_IOINST_net, 
        Y_DDR_DQ12_OUT_IOINST_net, D_DDR_DQ11_OUT_IOINST_net, 
        E_DDR_DQ11_OUT_IOINST_net, Y_DDR_DQ11_OUT_IOINST_net, 
        D_DDR_DQ10_OUT_IOINST_net, E_DDR_DQ10_OUT_IOINST_net, 
        Y_DDR_DQ10_OUT_IOINST_net, D_DDR_DQ9_OUT_IOINST_net, 
        E_DDR_DQ9_OUT_IOINST_net, Y_DDR_DQ9_OUT_IOINST_net, 
        D_DDR_DQ8_OUT_IOINST_net, E_DDR_DQ8_OUT_IOINST_net, 
        Y_DDR_DQ8_OUT_IOINST_net, D_DDR_DQ7_OUT_IOINST_net, 
        E_DDR_DQ7_OUT_IOINST_net, Y_DDR_DQ7_OUT_IOINST_net, 
        D_DDR_DQ6_OUT_IOINST_net, E_DDR_DQ6_OUT_IOINST_net, 
        Y_DDR_DQ6_OUT_IOINST_net, D_DDR_DQ5_OUT_IOINST_net, 
        E_DDR_DQ5_OUT_IOINST_net, Y_DDR_DQ5_OUT_IOINST_net, 
        D_DDR_DQ4_OUT_IOINST_net, E_DDR_DQ4_OUT_IOINST_net, 
        Y_DDR_DQ4_OUT_IOINST_net, D_DDR_DQ3_OUT_IOINST_net, 
        E_DDR_DQ3_OUT_IOINST_net, Y_DDR_DQ3_OUT_IOINST_net, 
        D_DDR_DQ2_OUT_IOINST_net, E_DDR_DQ2_OUT_IOINST_net, 
        Y_DDR_DQ2_OUT_IOINST_net, D_DDR_DQ1_OUT_IOINST_net, 
        E_DDR_DQ1_OUT_IOINST_net, Y_DDR_DQ1_OUT_IOINST_net, 
        D_DDR_DQ0_OUT_IOINST_net, E_DDR_DQ0_OUT_IOINST_net, 
        Y_DDR_DQ0_OUT_IOINST_net, D_DDR_DQS1_OUT_IOINST_net, 
        E_DDR_DQS1_OUT_IOINST_net, Y_DDR_DQS1_OUT_IOINST_net, 
        D_DDR_DQS0_OUT_IOINST_net, E_DDR_DQS0_OUT_IOINST_net, 
        Y_DDR_DQS0_OUT_IOINST_net, D_DDR_DM1_OUT_IOINST_net, 
        D_DDR_DM0_OUT_IOINST_net, D_DDR_RAM_RST_N_IOINST_net, 
        D_DDR_ODT0_IOINST_net, D_DDR_CKE0_IOINST_net, 
        D_DDR_CS0_IOINST_net, D_DDR_CK0_IOINST_net, 
        D_DDR_A5_IOINST_net, D_DDR_A4_IOINST_net, D_DDR_A3_IOINST_net, 
        D_DDR_A2_IOINST_net, D_DDR_A1_IOINST_net, D_DDR_A0_IOINST_net;
    assign FIC_3_APB_M_PADDR[31] = GND_net;
    assign FIC_3_APB_M_PADDR[29] = GND_net;
    
    BIBUF MSSIO9_OUT_IOINST (.D(D_MSSIO9_OUT_IOINST_net), .E(
        E_MSSIO9_OUT_IOINST_net), .Y(Y_MSSIO9_OUT_IOINST_net), .PAD(
        EMMC_DATA5_SD_VOLT_SEL));
    BIBUF MSSIO23_OUT_IOINST (.D(D_MSSIO23_OUT_IOINST_net), .E(
        E_MSSIO23_OUT_IOINST_net), .Y(Y_MSSIO23_OUT_IOINST_net), .PAD(
        USB_DATA5));
    OUTBUF DDR_CKE0_IOINST (.D(D_DDR_CKE0_IOINST_net), .PAD(CKE));
    OUTBUF DDR_CS0_IOINST (.D(D_DDR_CS0_IOINST_net), .PAD(CS));
    INBUF MSSIO14_IN_IOINST (.PAD(USB_CLK), .Y(Y_MSSIO14_IN_IOINST_net)
        );
    INV I_MSS_I2C_0_SDA_OE_M2F_INV (.A(I2C_0_SDA_OE_M2F_I_MSS_net), .Y(
        I2C_0_SDA_OE_M2F));
    INBUF MSSIO16_IN_IOINST (.PAD(USB_NXT), .Y(Y_MSSIO16_IN_IOINST_net)
        );
    OUTBUF MSSIO28_OUT_IOINST (.D(D_MSSIO28_OUT_IOINST_net), .PAD(
        MAC_1_MDC));
    OUTBUF MSSIO7_OUT_IOINST (.D(D_MSSIO7_OUT_IOINST_net), .PAD(
        EMMC_RSTN_SD_WP));
    INBUF_DIFF SGMII_RX1_IOINST (.PADP(SGMII_RX1_P), .PADN(SGMII_RX1_N)
        , .Y(Y_SGMII_RX1_IOINST_net));
    BIBUF DDR_DQ2_OUT_IOINST (.D(D_DDR_DQ2_OUT_IOINST_net), .E(
        E_DDR_DQ2_OUT_IOINST_net), .Y(Y_DDR_DQ2_OUT_IOINST_net), .PAD(
        DQ[2]));
    OUTBUF MSSIO12_OUT_IOINST (.D(D_MSSIO12_OUT_IOINST_net), .PAD(
        EMMC_UNUSED_SD_VOLT_DIR_0));
    INBUF MSSIO6_IN_IOINST (.PAD(EMMC_STRB_SD_CD), .Y(
        Y_MSSIO6_IN_IOINST_net));
    OUTBUF DDR_A4_IOINST (.D(D_DDR_A4_IOINST_net), .PAD(CA[4]));
    BIBUF MSSIO20_OUT_IOINST (.D(D_MSSIO20_OUT_IOINST_net), .E(
        E_MSSIO20_OUT_IOINST_net), .Y(Y_MSSIO20_OUT_IOINST_net), .PAD(
        USB_DATA2));
    BIBUF DDR_DQ3_OUT_IOINST (.D(D_DDR_DQ3_OUT_IOINST_net), .E(
        E_DDR_DQ3_OUT_IOINST_net), .Y(Y_DDR_DQ3_OUT_IOINST_net), .PAD(
        DQ[3]));
    OUTBUF DDR_DM0_OUT_IOINST (.D(D_DDR_DM0_OUT_IOINST_net), .PAD(
        DM[0]));
    OUTBUF MSSIO0_OUT_IOINST (.D(D_MSSIO0_OUT_IOINST_net), .PAD(
        EMMC_CLK_SD_CLK));
    OUTBUF DDR_A5_IOINST (.D(D_DDR_A5_IOINST_net), .PAD(CA[5]));
    OUTBUF DDR_DM1_OUT_IOINST (.D(D_DDR_DM1_OUT_IOINST_net), .PAD(
        DM[1]));
    OUTBUF DDR_A2_IOINST (.D(D_DDR_A2_IOINST_net), .PAD(CA[2]));
    BIBUF MSSIO32_OUT_IOINST (.D(D_MSSIO32_OUT_IOINST_net), .E(
        E_MSSIO32_OUT_IOINST_net), .Y(Y_MSSIO32_OUT_IOINST_net), .PAD(
        QSPI_DATA0));
    OUTBUF MSSIO36_OUT_IOINST (.D(D_MSSIO36_OUT_IOINST_net), .PAD(
        CAN_1_TX_EBL_N));
    BIBUF DDR_DQ4_OUT_IOINST (.D(D_DDR_DQ4_OUT_IOINST_net), .E(
        E_DDR_DQ4_OUT_IOINST_net), .Y(Y_DDR_DQ4_OUT_IOINST_net), .PAD(
        DQ[4]));
    OUTBUF DDR_ODT0_IOINST (.D(D_DDR_ODT0_IOINST_net), .PAD(ODT));
    BIBUF DDR_DQ9_OUT_IOINST (.D(D_DDR_DQ9_OUT_IOINST_net), .E(
        E_DDR_DQ9_OUT_IOINST_net), .Y(Y_DDR_DQ9_OUT_IOINST_net), .PAD(
        DQ[9]));
    BIBUF MSSIO29_OUT_IOINST (.D(D_MSSIO29_OUT_IOINST_net), .E(
        E_MSSIO29_OUT_IOINST_net), .Y(Y_MSSIO29_OUT_IOINST_net), .PAD(
        MAC_1_MDIO));
    OUTBUF MSSIO13_OUT_IOINST (.D(D_MSSIO13_OUT_IOINST_net), .PAD(
        EMMC_UNUSED_SD_VOLT_DIR_1_3));
    OUTBUF DDR_A1_IOINST (.D(D_DDR_A1_IOINST_net), .PAD(CA[1]));
    OUTBUF_DIFF SGMII_TX1_IOINST (.D(D_SGMII_TX1_IOINST_net), .PADP(
        SGMII_TX1_P), .PADN(SGMII_TX1_N));
    OUTBUF DDR_RAM_RST_N_IOINST (.D(D_DDR_RAM_RST_N_IOINST_net), .PAD(
        RESET_N));
    BIBUF MSSIO5_OUT_IOINST (.D(D_MSSIO5_OUT_IOINST_net), .E(
        E_MSSIO5_OUT_IOINST_net), .Y(Y_MSSIO5_OUT_IOINST_net), .PAD(
        EMMC_DATA3_SD_DATA3));
    BIBUF MSSIO33_OUT_IOINST (.D(D_MSSIO33_OUT_IOINST_net), .E(
        E_MSSIO33_OUT_IOINST_net), .Y(Y_MSSIO33_OUT_IOINST_net), .PAD(
        QSPI_DATA1));
    BIBUF MSSIO24_OUT_IOINST (.D(D_MSSIO24_OUT_IOINST_net), .E(
        E_MSSIO24_OUT_IOINST_net), .Y(Y_MSSIO24_OUT_IOINST_net), .PAD(
        USB_DATA6));
    BIBUF MSSIO18_OUT_IOINST (.D(D_MSSIO18_OUT_IOINST_net), .E(
        E_MSSIO18_OUT_IOINST_net), .Y(Y_MSSIO18_OUT_IOINST_net), .PAD(
        USB_DATA0));
    INBUF MSSIO15_IN_IOINST (.PAD(USB_DIR), .Y(Y_MSSIO15_IN_IOINST_net)
        );
    BIBUF MSSIO4_OUT_IOINST (.D(D_MSSIO4_OUT_IOINST_net), .E(
        E_MSSIO4_OUT_IOINST_net), .Y(Y_MSSIO4_OUT_IOINST_net), .PAD(
        EMMC_DATA2_SD_DATA2));
    OUTBUF_DIFF DDR_CK0_IOINST (.D(D_DDR_CK0_IOINST_net), .PADP(CK), 
        .PADN(CK_N));
    BIBUF MSSIO2_OUT_IOINST (.D(D_MSSIO2_OUT_IOINST_net), .E(
        E_MSSIO2_OUT_IOINST_net), .Y(Y_MSSIO2_OUT_IOINST_net), .PAD(
        EMMC_DATA0_SD_DATA0));
    BIBUF MSSIO27_OUT_IOINST (.D(D_MSSIO27_OUT_IOINST_net), .E(
        E_MSSIO27_OUT_IOINST_net), .Y(Y_MSSIO27_OUT_IOINST_net), .PAD(
        I2C_1_SDA));
    BIBUF_DIFF DDR_DQS0_OUT_IOINST (.Y(Y_DDR_DQS0_OUT_IOINST_net), .D(
        D_DDR_DQS0_OUT_IOINST_net), .E(E_DDR_DQS0_OUT_IOINST_net), 
        .PADP(DQS[0]), .PADN(DQS_N[0]));
    BIBUF MSSIO21_OUT_IOINST (.D(D_MSSIO21_OUT_IOINST_net), .E(
        E_MSSIO21_OUT_IOINST_net), .Y(Y_MSSIO21_OUT_IOINST_net), .PAD(
        USB_DATA3));
    BIBUF DDR_DQ14_OUT_IOINST (.D(D_DDR_DQ14_OUT_IOINST_net), .E(
        E_DDR_DQ14_OUT_IOINST_net), .Y(Y_DDR_DQ14_OUT_IOINST_net), 
        .PAD(DQ[14]));
    BIBUF DDR_DQ10_OUT_IOINST (.D(D_DDR_DQ10_OUT_IOINST_net), .E(
        E_DDR_DQ10_OUT_IOINST_net), .Y(Y_DDR_DQ10_OUT_IOINST_net), 
        .PAD(DQ[10]));
    INV I_MSS_I2C_0_SCL_OE_M2F_INV (.A(I2C_0_SCL_OE_M2F_I_MSS_net), .Y(
        I2C_0_SCL_OE_M2F));
    BIBUF MSSIO10_OUT_IOINST (.D(D_MSSIO10_OUT_IOINST_net), .E(
        E_MSSIO10_OUT_IOINST_net), .Y(Y_MSSIO10_OUT_IOINST_net), .PAD(
        EMMC_DATA6_SD_VOLT_EN));
    BIBUF DDR_DQ13_OUT_IOINST (.D(D_DDR_DQ13_OUT_IOINST_net), .E(
        E_DDR_DQ13_OUT_IOINST_net), .Y(Y_DDR_DQ13_OUT_IOINST_net), 
        .PAD(DQ[13]));
    BIBUF_DIFF DDR_DQS1_OUT_IOINST (.Y(Y_DDR_DQS1_OUT_IOINST_net), .D(
        D_DDR_DQS1_OUT_IOINST_net), .E(E_DDR_DQS1_OUT_IOINST_net), 
        .PADP(DQS[1]), .PADN(DQS_N[1]));
    BIBUF DDR_DQ11_OUT_IOINST (.D(D_DDR_DQ11_OUT_IOINST_net), .E(
        E_DDR_DQ11_OUT_IOINST_net), .Y(Y_DDR_DQ11_OUT_IOINST_net), 
        .PAD(DQ[11]));
    OUTBUF MSSIO30_OUT_IOINST (.D(D_MSSIO30_OUT_IOINST_net), .PAD(
        QSPI_CLK));
    OUTBUF DDR_A0_IOINST (.D(D_DDR_A0_IOINST_net), .PAD(CA[0]));
    INBUF_DIFF SGMII_RX0_IOINST (.PADP(SGMII_RX0_P), .PADN(SGMII_RX0_N)
        , .Y(Y_SGMII_RX0_IOINST_net));
    VCC VCC_inst (.Y(FIC_3_APB_M_PADDR[30]));
    BIBUF MSSIO8_OUT_IOINST (.D(D_MSSIO8_OUT_IOINST_net), .E(
        E_MSSIO8_OUT_IOINST_net), .Y(Y_MSSIO8_OUT_IOINST_net), .PAD(
        EMMC_DATA4_SD_POW));
    BIBUF DDR_DQ15_OUT_IOINST (.D(D_DDR_DQ15_OUT_IOINST_net), .E(
        E_DDR_DQ15_OUT_IOINST_net), .Y(Y_DDR_DQ15_OUT_IOINST_net), 
        .PAD(DQ[15]));
    OUTBUF_DIFF SGMII_TX0_IOINST (.D(D_SGMII_TX0_IOINST_net), .PADP(
        SGMII_TX0_P), .PADN(SGMII_TX0_N));
    BIBUF MSSIO19_OUT_IOINST (.D(D_MSSIO19_OUT_IOINST_net), .E(
        E_MSSIO19_OUT_IOINST_net), .Y(Y_MSSIO19_OUT_IOINST_net), .PAD(
        USB_DATA1));
    BIBUF DDR_DQ7_OUT_IOINST (.D(D_DDR_DQ7_OUT_IOINST_net), .E(
        E_DDR_DQ7_OUT_IOINST_net), .Y(Y_DDR_DQ7_OUT_IOINST_net), .PAD(
        DQ[7]));
    INBUF MSSIO35_IN_IOINST (.PAD(CAN_1_RXBUS), .Y(
        Y_MSSIO35_IN_IOINST_net));
    INBUF_DIFF REFCLK_IOINST (.PADP(REFCLK), .PADN(REFCLK_N), .Y(
        Y_REFCLK_IOINST_net));
    BIBUF MSSIO22_OUT_IOINST (.D(D_MSSIO22_OUT_IOINST_net), .E(
        E_MSSIO22_OUT_IOINST_net), .Y(Y_MSSIO22_OUT_IOINST_net), .PAD(
        USB_DATA4));
    GND GND_inst (.Y(GND_net));
    BIBUF DDR_DQ5_OUT_IOINST (.D(D_DDR_DQ5_OUT_IOINST_net), .E(
        E_DDR_DQ5_OUT_IOINST_net), .Y(Y_DDR_DQ5_OUT_IOINST_net), .PAD(
        DQ[5]));
    OUTBUF DDR_A3_IOINST (.D(D_DDR_A3_IOINST_net), .PAD(CA[3]));
    BIBUF MSSIO1_OUT_IOINST (.D(D_MSSIO1_OUT_IOINST_net), .E(
        E_MSSIO1_OUT_IOINST_net), .Y(Y_MSSIO1_OUT_IOINST_net), .PAD(
        EMMC_CMD_SD_CMD));
    MSS #( .MSS_CLK_DIV(1), .MSS_AHB_APB_CLK_DIV(4), .MSS_AXI_CLK_DIV(2)
        , .MSS_CLK_FREQ(600.0), .MSS_DDR_CLK_FREQ(800.0), .PROGRAM_NAME("pfsoc_mss")
        , .CORE_NAME("pfsoc_mss%2025.2"), .DIE("MPFS095T"), .PKG("FCSG325")
        , .BANK2_VDDI("3.3"), .BANK4_VDDI("1.8"), .BANK5_VDDI("3.3"), .DDR_SDRAM_TYPE("LPDDR4")
        , .REFCLK_IOSTD("LVDS25"), .SGMII_IOSTD("LVDS33"), .SGMII_RX0_IOSTD("LVDS33")
        , .SGMII_RX1_IOSTD("LVDS33"), .SGMII_TX0_IOSTD("LVDS33"), .SGMII_TX1_IOSTD("LVDS33")
        , .SPI0_CONTROL1_CFG_MODE(2'h0), .SPI1_CONTROL1_CFG_MODE(2'h0)
        , .DDR_SEGS_SEG0_0_ADDRESS_OFFSET(15'h7F80), .DDR_SEGS_SEG0_1_ADDRESS_OFFSET(15'h7030)
        , .DDR_SEGS_SEG1_2_ADDRESS_OFFSET(15'h7FB0), .DDR_SEGS_SEG1_3_ADDRESS_OFFSET(15'h0)
        , .DDR_SEGS_SEG1_4_ADDRESS_OFFSET(15'h7FA0), .DDR_SEGS_SEG1_5_ADDRESS_OFFSET(15'h0)
        , .DDR_SEGS_SEG1_6_ADDRESS_OFFSET(15'h0), .DDR_DDRC_CFG_AXI_START_ADDRESS_AXI1_0(32'h0)
        , .DDR_DDRC_CFG_AXI_START_ADDRESS_AXI1_1(32'h0), .DDR_DDRC_CFG_AXI_START_ADDRESS_AXI2_0(32'h0)
        , .DDR_DDRC_CFG_AXI_START_ADDRESS_AXI2_1(32'h0), .DDR_DDRC_CFG_AXI_END_ADDRESS_AXI1_0(32'hFFFFFFFF)
        , .DDR_DDRC_CFG_AXI_END_ADDRESS_AXI1_1(32'h3), .DDR_DDRC_CFG_AXI_END_ADDRESS_AXI2_0(32'hFFFFFFFF)
        , .DDR_DDRC_CFG_AXI_END_ADDRESS_AXI2_1(32'h3), .DDR_DDRC_CFG_MEM_START_ADDRESS_AXI1_0(32'h0)
        , .DDR_DDRC_CFG_MEM_START_ADDRESS_AXI1_1(32'h0), .DDR_DDRC_CFG_MEM_START_ADDRESS_AXI2_0(32'h0)
        , .DDR_DDRC_CFG_MEM_START_ADDRESS_AXI2_1(32'h0), .MSSIO_IOMUX0_CR_SPI0_FABRIC(1'h1)
        , .MSSIO_IOMUX0_CR_SPI1_FABRIC(1'h0), .MSSIO_IOMUX0_CR_I2C0_FABRIC(1'h1)
        , .MSSIO_IOMUX0_CR_I2C1_FABRIC(1'h0), .MSSIO_IOMUX0_CR_CAN0_FABRIC(1'h1)
        , .MSSIO_IOMUX0_CR_CAN1_FABRIC(1'h0), .MSSIO_IOMUX0_CR_QSPI_FABRIC(1'h0)
        , .MSSIO_IOMUX0_CR_MMUART0_FABRIC(1'h1), .MSSIO_IOMUX0_CR_MMUART1_FABRIC(1'h1)
        , .MSSIO_IOMUX0_CR_MMUART2_FABRIC(1'h1), .MSSIO_IOMUX0_CR_MMUART3_FABRIC(1'h1)
        , .MSSIO_IOMUX0_CR_MMUART4_FABRIC(1'h1), .MSSIO_IOMUX0_CR_MDIO0_FABRIC(1'h0)
        , .MSSIO_IOMUX0_CR_MDIO1_FABRIC(1'h0), .MSSIO_IOMUX1_CR_PAD0(4'h1)
        , .MSSIO_IOMUX1_CR_PAD1(4'h1), .MSSIO_IOMUX1_CR_PAD2(4'h1), .MSSIO_IOMUX1_CR_PAD3(4'h1)
        , .MSSIO_IOMUX1_CR_PAD4(4'h1), .MSSIO_IOMUX1_CR_PAD5(4'h1), .MSSIO_IOMUX1_CR_PAD6(4'h1)
        , .MSSIO_IOMUX1_CR_PAD7(4'h1), .MSSIO_IOMUX2_CR_PAD8(4'h1), .MSSIO_IOMUX2_CR_PAD9(4'h1)
        , .MSSIO_IOMUX2_CR_PAD10(4'h1), .MSSIO_IOMUX2_CR_PAD11(4'h1), .MSSIO_IOMUX2_CR_PAD12(4'hF)
        , .MSSIO_IOMUX2_CR_PAD13(4'hF), .MSSIO_IOMUX3_CR_PAD14(4'h4), .MSSIO_IOMUX3_CR_PAD15(4'h4)
        , .MSSIO_IOMUX3_CR_PAD16(4'h4), .MSSIO_IOMUX3_CR_PAD17(4'h4), .MSSIO_IOMUX3_CR_PAD18(4'h4)
        , .MSSIO_IOMUX3_CR_PAD19(4'h4), .MSSIO_IOMUX3_CR_PAD20(4'h4), .MSSIO_IOMUX3_CR_PAD21(4'h4)
        , .MSSIO_IOMUX4_CR_PAD22(4'h4), .MSSIO_IOMUX4_CR_PAD23(4'h4), .MSSIO_IOMUX4_CR_PAD24(4'h4)
        , .MSSIO_IOMUX4_CR_PAD25(4'h4), .MSSIO_IOMUX4_CR_PAD26(4'h6), .MSSIO_IOMUX4_CR_PAD27(4'h6)
        , .MSSIO_IOMUX4_CR_PAD28(4'h8), .MSSIO_IOMUX4_CR_PAD29(4'h8), .MSSIO_IOMUX5_CR_PAD30(4'h2)
        , .MSSIO_IOMUX5_CR_PAD31(4'h2), .MSSIO_IOMUX5_CR_PAD32(4'h2), .MSSIO_IOMUX5_CR_PAD33(4'h2)
        , .MSSIO_IOMUX5_CR_PAD34(4'h7), .MSSIO_IOMUX5_CR_PAD35(4'h7), .MSSIO_IOMUX5_CR_PAD36(4'h7)
        , .MSSIO_IOMUX5_CR_PAD37(4'hF), .MSSIO_IOMUX6_CR_VLT_SEL(1'h0)
        , .MSSIO_IOMUX6_CR_VLT_EN(1'h0), .MSSIO_IOMUX6_CR_VLT_CMD_DIR(1'h0)
        , .MSSIO_IOMUX6_CR_VLT_DIR_0(1'h0), .MSSIO_IOMUX6_CR_VLT_DIR_1_3(1'h0)
        , .MSSIO_IOMUX6_CR_SD_LED(1'h0), .MSSIO_IOMUX6_CR_SD_VOLT_0(1'h0)
        , .MSSIO_IOMUX6_CR_SD_VOLT_1(1'h0), .MSSIO_IOMUX6_CR_SD_VOLT_2(1'h0)
        , .MSSIO_MSSIO_BANK2_CFG_CR_BANK_PCODE(6'h7), .MSSIO_MSSIO_BANK2_CFG_CR_BANK_NCODE(6'h9)
        , .MSSIO_MSSIO_BANK2_CFG_CR_VS(4'h8), .MSSIO_MSSIO_BANK4_CFG_CR_BANK_PCODE(6'hD)
        , .MSSIO_MSSIO_BANK4_CFG_CR_BANK_NCODE(6'hA), .MSSIO_MSSIO_BANK4_CFG_CR_VS(4'h4)
        , .SGMII_SGMII_MODE_REG_BC_VS(4'h8), .SGMII_SGMII_MODE_REG_PLL_EN(1'h1)
        , .SGMII_SGMII_MODE_REG_DLL_EN(1'h1), .SGMII_DYN_CNTL_REG_PLL_SOFT_RESET_PERIPH(1'h0)
        , .SGMII_DYN_CNTL_REG_DLL_SOFT_RESET_PERIPH(1'h0), .SGMII_DYN_CNTL_REG_PVT_SOFT_RESET_PERIPH(1'h0)
        , .SGMII_DYN_CNTL_REG_BC_SOFT_RESET_PERIPH(1'h0), .SGMII_SGMII_MODE_REG_TX0_EN(1'h1)
        , .SGMII_SGMII_MODE_REG_RX0_EN(1'h1), .SGMII_SGMII_MODE_REG_CH0_CDR_RESET_B(1'h1)
        , .SGMII_DYN_CNTL_REG_LANE0_SOFT_RESET_PERIPH(1'h0), .SGMII_CH0_CNTL_REG_TX0_WPU_P(1'h0)
        , .SGMII_CH0_CNTL_REG_TX0_WPD_P(1'h0), .SGMII_CH0_CNTL_REG_TX0_SLEW_P(2'h0)
        , .SGMII_CH0_CNTL_REG_TX0_DRV_P(4'h7), .SGMII_CH0_CNTL_REG_TX0_ODT_P(4'h7)
        , .SGMII_CH0_CNTL_REG_TX0_ODT_STATIC_P(3'h7), .SGMII_CH0_CNTL_REG_RX0_WPU_P(1'h0)
        , .SGMII_CH0_CNTL_REG_RX0_WPD_P(1'h0), .SGMII_CH0_CNTL_REG_RX0_IBUFMD_P(3'h4)
        , .SGMII_CH0_CNTL_REG_RX0_ODT_P(4'h7), .SGMII_CH0_CNTL_REG_RX0_ODT_STATIC_P(3'h3)
        , .SGMII_SGMII_MODE_REG_TX1_EN(1'h1), .SGMII_SGMII_MODE_REG_RX1_EN(1'h1)
        , .SGMII_SGMII_MODE_REG_CH1_CDR_RESET_B(1'h1), .SGMII_DYN_CNTL_REG_LANE1_SOFT_RESET_PERIPH(1'h0)
        , .SGMII_CH1_CNTL_REG_TX1_WPU_P(1'h0), .SGMII_CH1_CNTL_REG_TX1_WPD_P(1'h0)
        , .SGMII_CH1_CNTL_REG_TX1_SLEW_P(2'h0), .SGMII_CH1_CNTL_REG_TX1_DRV_P(4'h7)
        , .SGMII_CH1_CNTL_REG_TX1_ODT_P(4'h7), .SGMII_CH1_CNTL_REG_TX1_ODT_STATIC_P(3'h7)
        , .SGMII_CH1_CNTL_REG_RX1_WPU_P(1'h0), .SGMII_CH1_CNTL_REG_RX1_WPD_P(1'h0)
        , .SGMII_CH1_CNTL_REG_RX1_IBUFMD_P(3'h4), .SGMII_CH1_CNTL_REG_RX1_ODT_P(4'h7)
        , .SGMII_CH1_CNTL_REG_RX1_ODT_STATIC_P(3'h3), .SGMII_SGMII_MODE_REG_PVT_EN(1'h1)
        , .SGMII_SGMII_MODE_REG_BC_VRGEN_EN(1'h1), .SGMII_RECAL_CNTL_REG_PVT_CALIB_START(1'h1)
        , .SGMII_RECAL_CNTL_REG_PVT_CALIB_LOCK(1'h1), .SGMII_DYN_CNTL_REG_CLKMUX_SOFT_RESET_PERIPH(1'h0)
        , .SGMII_CLK_CNTL_REG_REFCLK_EN_RXMODE_P(2'h3), .SGMII_CLK_CNTL_REG_REFCLK_EN_RXMODE_N(2'h3)
        , .CLK_SGMII_CFM_CLK_XCVR_EN_RXMODE_P(2'h3), .CLK_SGMII_CFM_CLK_XCVR_EN_RXMODE_N(2'h3)
        , .SGMII_SGMII_MODE_REG_REFCLK_EN_UDRIVE_P(1'h0), .SGMII_SGMII_MODE_REG_REFCLK_EN_UDRIVE_N(1'h0)
        , .CLK_SGMII_CFM_CLK_XCVR_EN_UDRIVE_P(1'h0), .CLK_SGMII_CFM_CLK_XCVR_EN_UDRIVE_N(1'h0)
        , .SGMII_SGMII_MODE_REG_REFCLK_EN_RDIFF(1'h1), .CLK_SGMII_CFM_CLK_XCVR_EN_RDIFF(1'h1)
        , .SGMII_CLK_CNTL_REG_REFCLK_EN_TERM_P(2'h0), .SGMII_CLK_CNTL_REG_REFCLK_EN_TERM_N(2'h0)
        , .CLK_SGMII_CFM_CLK_XCVR_EN_TERM_P(2'h0), .CLK_SGMII_CFM_CLK_XCVR_EN_TERM_N(2'h0)
        , .SGMII_SGMII_MODE_REG_REFCLK_EN_INS_HYST_P(1'h0), .SGMII_SGMII_MODE_REG_REFCLK_EN_INS_HYST_N(1'h0)
        , .CLK_SGMII_CFM_CLK_XCVR_EN_INS_HYST_P(1'h0), .CLK_SGMII_CFM_CLK_XCVR_EN_INS_HYST_N(1'h0)
        , .SGMII_CLK_CNTL_REG_REFCLK_CLKBUF_EN_PULLUP(1'h0), .CLK_SGMII_CFM_CLK_XCVR_CLKBUF_EN_PULLUP(1'h0)
        , .MSSIO_MSSIO_BANK4_IO_CFG_0_1_CR_IO_CFG_0(16'h0928), .MSSIO_MSSIO_BANK4_IO_CFG_0_1_CR_IO_CFG_1(16'h0928)
        , .MSSIO_MSSIO_BANK4_IO_CFG_2_3_CR_IO_CFG_2(16'h0928), .MSSIO_MSSIO_BANK4_IO_CFG_2_3_CR_IO_CFG_3(16'h0928)
        , .MSSIO_MSSIO_BANK4_IO_CFG_4_5_CR_IO_CFG_4(16'h0928), .MSSIO_MSSIO_BANK4_IO_CFG_4_5_CR_IO_CFG_5(16'h0928)
        , .MSSIO_MSSIO_BANK4_IO_CFG_6_7_CR_IO_CFG_6(16'h0928), .MSSIO_MSSIO_BANK4_IO_CFG_6_7_CR_IO_CFG_7(16'h0928)
        , .MSSIO_MSSIO_BANK4_IO_CFG_8_9_CR_IO_CFG_8(16'h0928), .MSSIO_MSSIO_BANK4_IO_CFG_8_9_CR_IO_CFG_9(16'h0928)
        , .MSSIO_MSSIO_BANK4_IO_CFG_10_11_CR_IO_CFG_10(16'h0928), .MSSIO_MSSIO_BANK4_IO_CFG_10_11_CR_IO_CFG_11(16'h0928)
        , .MSSIO_MSSIO_BANK4_IO_CFG_12_13_CR_IO_CFG_12(16'h0928), .MSSIO_MSSIO_BANK4_IO_CFG_12_13_CR_IO_CFG_13(16'h0928)
        , .MSSIO_MSSIO_BANK2_IO_CFG_0_1_CR_IO_CFG_0(16'h0829), .MSSIO_MSSIO_BANK2_IO_CFG_0_1_CR_IO_CFG_1(16'h0829)
        , .MSSIO_MSSIO_BANK2_IO_CFG_2_3_CR_IO_CFG_2(16'h0829), .MSSIO_MSSIO_BANK2_IO_CFG_2_3_CR_IO_CFG_3(16'h0829)
        , .MSSIO_MSSIO_BANK2_IO_CFG_4_5_CR_IO_CFG_4(16'h0829), .MSSIO_MSSIO_BANK2_IO_CFG_4_5_CR_IO_CFG_5(16'h0829)
        , .MSSIO_MSSIO_BANK2_IO_CFG_6_7_CR_IO_CFG_6(16'h0829), .MSSIO_MSSIO_BANK2_IO_CFG_6_7_CR_IO_CFG_7(16'h0829)
        , .MSSIO_MSSIO_BANK2_IO_CFG_8_9_CR_IO_CFG_8(16'h0829), .MSSIO_MSSIO_BANK2_IO_CFG_8_9_CR_IO_CFG_9(16'h0829)
        , .MSSIO_MSSIO_BANK2_IO_CFG_10_11_CR_IO_CFG_10(16'h0829), .MSSIO_MSSIO_BANK2_IO_CFG_10_11_CR_IO_CFG_11(16'h0829)
        , .MSSIO_MSSIO_BANK2_IO_CFG_12_13_CR_IO_CFG_12(16'h0829), .MSSIO_MSSIO_BANK2_IO_CFG_12_13_CR_IO_CFG_13(16'h0829)
        , .MSSIO_MSSIO_BANK2_IO_CFG_14_15_CR_IO_CFG_14(16'h0829), .MSSIO_MSSIO_BANK2_IO_CFG_14_15_CR_IO_CFG_15(16'h0829)
        , .MSSIO_MSSIO_BANK2_IO_CFG_16_17_CR_IO_CFG_16(16'h0829), .MSSIO_MSSIO_BANK2_IO_CFG_16_17_CR_IO_CFG_17(16'h0829)
        , .MSSIO_MSSIO_BANK2_IO_CFG_18_19_CR_IO_CFG_18(16'h0829), .MSSIO_MSSIO_BANK2_IO_CFG_18_19_CR_IO_CFG_19(16'h0829)
        , .MSSIO_MSSIO_BANK2_IO_CFG_20_21_CR_IO_CFG_20(16'h0829), .MSSIO_MSSIO_BANK2_IO_CFG_20_21_CR_IO_CFG_21(16'h0829)
        , .MSSIO_MSSIO_BANK2_IO_CFG_22_23_CR_IO_CFG_22(16'h0829), .MSSIO_MSSIO_BANK2_IO_CFG_22_23_CR_IO_CFG_23(16'h0829)
        , .GENERAL_GPIO_CR_GPIO0_SOFT_RESET_SELECT(2'h3), .GENERAL_GPIO_CR_GPIO1_SOFT_RESET_SELECT(3'h7)
        , .GENERAL_GPIO_CR_GPIO2_SOFT_RESET_SELECT(4'hF), .GENERAL_CRYPTO_CR_INFO_MSS_MODE(2'h0)
        , .DDR_DDRC_CFG_CHIPADDR_MAP_CFG_CHIPADDR_MAP(32'h00001D), .DDR_DDRC_CFG_BANKADDR_MAP_0_CFG_BANKADDR_MAP_0(32'h00C2CA)
        , .DDR_DDRC_CFG_ROWADDR_MAP_0_CFG_ROWADDR_MAP_0(32'h9140F38D)
        , .DDR_DDRC_CFG_ROWADDR_MAP_1_CFG_ROWADDR_MAP_1(32'h75955134)
        , .DDR_DDRC_CFG_ROWADDR_MAP_2_CFG_ROWADDR_MAP_2(32'h71B69961)
        , .DDR_DDRC_CFG_ROWADDR_MAP_3_CFG_ROWADDR_MAP_3(32'h000), .DDR_DDRC_CFG_COLADDR_MAP_0_CFG_COLADDR_MAP_0(32'h440C2040)
        , .DDR_DDRC_CFG_COLADDR_MAP_1_CFG_COLADDR_MAP_1(32'h02481C61)
        , .DDR_DDRC_CFG_COLADDR_MAP_2_CFG_COLADDR_MAP_2(32'h00000000)
        , .DDR_DDRC_CFG_MEM_COLBITS_CFG_MEM_COLBITS(32'hA), .DDR_DDRC_CFG_MEM_ROWBITS_CFG_MEM_ROWBITS(32'h10)
        , .DDR_DDRC_CFG_MEM_BANKBITS_CFG_MEM_BANKBITS(32'h3), .DDR_DDRC_CFG_CL_CFG_CL(32'h5)
        , .DDR_DDRC_CFG_CWL_CFG_CWL(32'h5), .DDR_DDRC_CFG_NUM_RANKS_CFG_NUM_RANKS(32'h1)
        , .DDR_DDRC_CFG_ZQINIT_CAL_DURATION_CFG_ZQINIT_CAL_DURATION(32'h0)
        , .DDR_DDRC_CFG_ZQ_CAL_L_DURATION_CFG_ZQ_CAL_L_DURATION(32'h0)
        , .DDR_DDRC_CFG_ZQ_CAL_S_DURATION_CFG_ZQ_CAL_S_DURATION(32'h0)
        , .DDR_DDRC_CFG_ODT_RD_MAP_CS0_CFG_ODT_RD_MAP_CS0(32'h0), .DDR_DDRC_CFG_ODT_RD_MAP_CS1_CFG_ODT_RD_MAP_CS1(32'h0)
        , .DDR_DDRC_CFG_ODT_WR_MAP_CS0_CFG_ODT_WR_MAP_CS0(32'h0), .DDR_DDRC_CFG_ODT_WR_MAP_CS1_CFG_ODT_WR_MAP_CS1(32'h0)
        , .DDR_DDRC_CFG_RAS_CFG_RAS(32'h22), .DDR_DDRC_CFG_RCD_CFG_RCD(32'hF)
        , .DDR_DDRC_CFG_RRD_CFG_RRD(32'h8), .DDR_DDRC_CFG_RP_CFG_RP(32'h11)
        , .DDR_DDRC_CFG_RC_CFG_RC(32'h33), .DDR_DDRC_CFG_FAW_CFG_FAW(32'h20)
        , .DDR_DDRC_CFG_RFC_CFG_RFC(32'h130), .DDR_DDRC_CFG_RTP_CFG_RTP(32'h8)
        , .DDR_DDRC_CFG_WR_CFG_WR(32'h10), .DDR_DDRC_CFG_REF_PER_CFG_REF_PER(32'hC34)
        , .DDR_DDRC_CFG_STARTUP_DELAY_CFG_STARTUP_DELAY(32'h27100), .DDR_DDRC_CFG_ZQ_CAL_PER_CFG_ZQ_CAL_PER(32'h27100)
        , .DDR_DDRC_CFG_WTR_CFG_WTR(32'h8), .DDR_DDRC_CFG_MOD_CFG_MOD(32'hC)
        , .DDR_DDRC_CFG_XS_CFG_XS(32'h5), .DDR_DDRC_CFG_XPR_CFG_XPR(32'h5)
        , .DDR_DDRC_CFG_MANUAL_ADDRESS_MAP_CFG_MANUAL_ADDRESS_MAP(32'h0)
        , .DDR_DDRC_CFG_LOOKAHEAD_PCH_CFG_LOOKAHEAD_PCH(32'h0), .DDR_DDRC_CFG_LOOKAHEAD_ACT_CFG_LOOKAHEAD_ACT(32'h0)
        , .DDR_DDRC_CFG_AUTO_REF_EN_CFG_AUTO_REF_EN(32'h1), .DDR_DDRC_PHY_PC_RANK_PHY_PC_RANK(32'h1)
        , .DDR_DDRC_PHY_RANKS_TO_TRAIN_PHY_RANKS_TO_TRAIN(32'h1), .DDR_DDRC_CFG_RMW_EN_CFG_RMW_EN(32'h1)
        , .DDR_DDRC_CFG_ECC_CORRECTION_EN_CFG_ECC_CORRECTION_EN(32'h0)
        , .DDR_DDRC_CFG_ONLY_SRANK_CMDS_CFG_ONLY_SRANK_CMDS(32'h0), .DDR_DDRC_INIT_RDIMM_COMPLETE_INIT_RDIMM_COMPLETE(32'h0)
        , .DDR_DDRC_CFG_DM_EN_CFG_DM_EN(32'h0), .DDR_DDRC_CFG_AL_MODE_CFG_AL_MODE(32'h0)
        , .DDR_DDRC_CFG_BL_MODE_CFG_BL_MODE(32'h0), .DDR_DDRC_CFG_RTT_WR_CFG_RTT_WR(32'h0)
        , .DDR_DDRC_CFG_SRT_CFG_SRT(32'h0), .DDR_DDRC_CFG_ADDR_MIRROR_CFG_ADDR_MIRROR(32'h0)
        , .DDR_DDRC_CFG_ZQ_CAL_TYPE_CFG_ZQ_CAL_TYPE(32'h1), .DDR_DDRC_CFG_REGDIMM_CFG_REGDIMM(32'h0)
        , .DDR_DDRC_CFG_PASR_CFG_PASR(32'h0), .DDR_DDRC_CFG_BT_CFG_BT(32'h0)
        , .DDR_DDRC_CFG_DS_CFG_DS(32'h6), .DDR_DDRC_CFG_RTT_CFG_RTT(32'h2)
        , .DDR_DDRC_CFG_BANKADDR_MAP_1_CFG_BANKADDR_MAP_1(32'h0), .DDR_DDRC_CFG_NIBBLE_DEVICES_CFG_NIBBLE_DEVICES(32'h0)
        , .DDR_DDRC_CTRLR_SOFT_RESET_N_CTRLR_SOFT_RESET_N(32'h1), .DDR_DDRC_CFG_READ_TO_WRITE_CFG_READ_TO_WRITE(32'hF)
        , .DDR_DDRC_CFG_WRITE_TO_WRITE_CFG_WRITE_TO_WRITE(32'hF), .DDR_DDRC_CFG_READ_TO_READ_CFG_READ_TO_READ(32'hF)
        , .DDR_DDRC_CFG_WRITE_TO_READ_CFG_WRITE_TO_READ(32'h1F), .DDR_DDRC_CFG_READ_TO_WRITE_ODT_CFG_READ_TO_WRITE_ODT(32'hF)
        , .DDR_DDRC_CFG_WRITE_TO_WRITE_ODT_CFG_WRITE_TO_WRITE_ODT(32'h0)
        , .DDR_DDRC_CFG_READ_TO_READ_ODT_CFG_READ_TO_READ_ODT(32'h1), .DDR_DDRC_CFG_WRITE_TO_READ_ODT_CFG_WRITE_TO_READ_ODT(32'h1)
        , .DDR_DDRC_CFG_MIN_READ_IDLE_CFG_MIN_READ_IDLE(32'h7), .DDR_DDRC_CFG_QOFF_CFG_QOFF(32'h0)
        , .DDR_DDRC_CFG_DLL_DISABLE_CFG_DLL_DISABLE(32'h0), .DDR_DDRC_CFG_ODT_RD_MAP_CS2_CFG_ODT_RD_MAP_CS2(32'h0)
        , .DDR_DDRC_CFG_ODT_RD_MAP_CS3_CFG_ODT_RD_MAP_CS3(32'h0), .DDR_DDRC_CFG_ODT_RD_MAP_CS4_CFG_ODT_RD_MAP_CS4(32'h0)
        , .DDR_DDRC_CFG_ODT_RD_MAP_CS5_CFG_ODT_RD_MAP_CS5(32'h0), .DDR_DDRC_CFG_ODT_RD_MAP_CS6_CFG_ODT_RD_MAP_CS6(32'h0)
        , .DDR_DDRC_CFG_ODT_RD_MAP_CS7_CFG_ODT_RD_MAP_CS7(32'h0), .DDR_DDRC_CFG_ODT_WR_MAP_CS2_CFG_ODT_WR_MAP_CS2(32'h0)
        , .DDR_DDRC_CFG_ODT_WR_MAP_CS3_CFG_ODT_WR_MAP_CS3(32'h0), .DDR_DDRC_CFG_ODT_WR_MAP_CS4_CFG_ODT_WR_MAP_CS4(32'h0)
        , .DDR_DDRC_CFG_ODT_WR_MAP_CS5_CFG_ODT_WR_MAP_CS5(32'h0), .DDR_DDRC_CFG_ODT_WR_MAP_CS6_CFG_ODT_WR_MAP_CS6(32'h0)
        , .DDR_DDRC_CFG_ODT_WR_MAP_CS7_CFG_ODT_WR_MAP_CS7(32'h0), .DDR_DDRC_CFG_ODT_RD_TURN_ON_CFG_ODT_RD_TURN_ON(32'h0)
        , .DDR_DDRC_CFG_ODT_WR_TURN_ON_CFG_ODT_WR_TURN_ON(32'h0), .DDR_DDRC_CFG_ODT_RD_TURN_OFF_CFG_ODT_RD_TURN_OFF(32'h0)
        , .DDR_DDRC_CFG_ODT_WR_TURN_OFF_CFG_ODT_WR_TURN_OFF(32'h0), .DDR_DDRC_CFG_EMR3_CFG_EMR3(32'h0)
        , .DDR_DDRC_CFG_TWO_T_CFG_TWO_T(32'h0), .DDR_DDRC_CFG_TWO_T_SEL_CYCLE_CFG_TWO_T_SEL_CYCLE(32'h1)
        , .DDR_DDRC_CFG_TDQS_CFG_TDQS(32'h0), .DDR_DDRC_CFG_AUTO_SR_CFG_AUTO_SR(32'h0)
        , .DDR_DDRC_CFG_AUTO_ZQ_CAL_EN_CFG_AUTO_ZQ_CAL_EN(32'h1), .DDR_DDRC_CFG_MEMORY_TYPE_CFG_MEMORY_TYPE(32'h400)
        , .DDR_DDRC_CFG_QUAD_RANK_CFG_QUAD_RANK(32'h0), .DDR_DDRC_CFG_EARLY_RANK_TO_WR_START_CFG_EARLY_RANK_TO_WR_START(32'h0)
        , .DDR_DDRC_CFG_EARLY_RANK_TO_RD_START_CFG_EARLY_RANK_TO_RD_START(32'h0)
        , .DDR_DDRC_CFG_CAL_READ_PERIOD_CFG_CAL_READ_PERIOD(32'h0), .DDR_DDRC_CFG_NUM_CAL_READS_CFG_NUM_CAL_READS(32'h1)
        , .DDR_DDRC_CFG_CTRLR_INIT_DISABLE_CFG_CTRLR_INIT_DISABLE(32'h0)
        , .DDR_DDRC_CFG_RDIMM_LAT_CFG_RDIMM_LAT(32'h0), .DDR_DDRC_CFG_CTRLUPD_TRIG_CFG_CTRLUPD_TRIG(32'h0)
        , .DDR_DDRC_CFG_CTRLUPD_START_DELAY_CFG_CTRLUPD_START_DELAY(32'h0)
        , .DDR_DDRC_CFG_DFI_T_CTRLUPD_MAX_CFG_DFI_T_CTRLUPD_MAX(32'h0)
        , .DDR_DDRC_CFG_DFI_T_RDDATA_EN_CFG_DFI_T_RDDATA_EN(32'h15), .DDR_DDRC_CFG_DFI_T_PHY_WRLAT_CFG_DFI_T_PHY_WRLAT(32'h3)
        , .DDR_DDRC_PHY_DFI_INIT_START_PHY_DFI_INIT_START(32'h1), .DDR_DDRC_PHY_RESET_CONTROL_PHY_RESET_CONTROL(32'h8001)
        , .DDR_DDRC_PHY_GATE_TRAIN_DELAY_PHY_GATE_TRAIN_DELAY(32'h3F)
        , .DDR_DDRC_PHY_EYE_TRAIN_DELAY_PHY_EYE_TRAIN_DELAY(32'h3F), .DDR_DDRC_PHY_TRAIN_STEP_ENABLE_PHY_TRAIN_STEP_ENABLE(32'h18)
        , .DDR_DDRC_PHY_INDPNDT_TRAINING_PHY_INDPNDT_TRAINING(32'h1), .DDR_DDRC_CFG_DQ_WIDTH_CFG_DQ_WIDTH(32'h1)
        , .DDR_DDRC_CFG_CA_PARITY_ERR_STATUS_CFG_CA_PARITY_ERR_STATUS(32'h0)
        , .DDR_DDRC_CFG_PARITY_RDIMM_DELAY_CFG_PARITY_RDIMM_DELAY(32'h0)
        , .DDR_DDRC_CFG_DFI_T_PHY_RDLAT_CFG_DFI_T_PHY_RDLAT(32'h6), .DDR_DDRC_CFG_DATA_MASK_CFG_DATA_MASK(32'h1)
        , .DDR_MODEL_DATA_LANES_USED_DATA_LANES(3'h2), .DDR_DDRC_CFG_CCD_S_CFG_CCD_S(32'h5)
        , .DDR_DDRC_CFG_CCD_L_CFG_CCD_L(32'h6), .DDR_DDRC_CFG_RRD_S_CFG_RRD_S(32'h4)
        , .DDR_DDRC_CFG_RRD_L_CFG_RRD_L(32'h3), .DDR_DDRC_CFG_WTR_S_CFG_WTR_S(32'h3)
        , .DDR_DDRC_CFG_WTR_L_CFG_WTR_L(32'h3), .DDR_DDRC_CFG_WTR_S_CRC_DM_CFG_WTR_S_CRC_DM(32'h3)
        , .DDR_DDRC_CFG_WTR_L_CRC_DM_CFG_WTR_L_CRC_DM(32'h3), .DDR_DDRC_CFG_WR_CRC_DM_CFG_WR_CRC_DM(32'h6)
        , .DDR_DDRC_CFG_VREFDQ_TRN_VALUE_CFG_VREFDQ_TRN_VALUE(32'h17)
        , .DDR_DDRC_CFG_RFC1_CFG_RFC1(32'h36), .DDR_DDRC_CFG_RFC2_CFG_RFC2(32'h36)
        , .DDR_DDRC_CFG_RFC4_CFG_RFC4(32'h36), .DDR_DDRC_CFG_FINE_GRAN_REF_MODE_CFG_FINE_GRAN_REF_MODE(32'h0)
        , .DDR_DDRC_CFG_RD_PREAMBLE_CFG_RD_PREAMBLE(32'h0), .DDR_DDRC_CFG_SR_ABORT_CFG_SR_ABORT(32'h0)
        , .DDR_DDRC_CFG_INT_VREF_MON_CFG_INT_VREF_MON(32'h0), .DDR_DDRC_CFG_TEMP_CTRL_REF_MODE_CFG_TEMP_CTRL_REF_MODE(32'h0)
        , .DDR_DDRC_CFG_TEMP_CTRL_REF_RANGE_CFG_TEMP_CTRL_REF_RANGE(32'h0)
        , .DDR_DDRC_CFG_RTT_PARK_CFG_RTT_PARK(32'h0), .DDR_DDRC_CFG_ODT_INBUF_4_PD_CFG_ODT_INBUF_4_PD(32'h0)
        , .DDR_DDRC_CFG_CA_PARITY_LATENCY_CFG_CA_PARITY_LATENCY(32'h0)
        , .DDR_DDRC_CFG_VREFDQ_TRN_ENABLE_CFG_VREFDQ_TRN_ENABLE(32'h1)
        , .DDR_DDRC_CFG_VREFDQ_TRN_RANGE_CFG_VREFDQ_TRN_RANGE(32'h1), .DDR_DDRC_CFG_LP_ASR_CFG_LP_ASR(32'h0)
        , .DDR_DDRC_CFG_WR_PREAMBLE_CFG_WR_PREAMBLE(32'h1), .DDR_DDRC_CFG_RFC_DLR1_CFG_RFC_DLR1(32'h48)
        , .DDR_DDRC_CFG_RFC_DLR2_CFG_RFC_DLR2(32'h2C), .DDR_DDRC_CFG_RFC_DLR4_CFG_RFC_DLR4(32'h20)
        , .DDR_DDRC_CFG_RRD_DLR_CFG_RRD_DLR(32'h4), .DDR_DDRC_CFG_FAW_DLR_CFG_FAW_DLR(32'h10)
        , .DDR_DDRC_CFG_BG_INTERLEAVE_CFG_BG_INTERLEAVE(32'h1), .DDR_DDRC_CFG_MRR_CFG_MRR(32'h8)
        , .DDR_DDRC_CFG_MRW_CFG_MRW(32'hA), .DDR_DDRC_CFG_XP_CFG_XP(32'h6)
        , .DDR_DDRC_CFG_XSR_CFG_XSR(32'h1F), .DDR_DDRC_CFG_INIT_DURATION_CFG_INIT_DURATION(32'h640)
        , .DDR_DDRC_CFG_ZQ_CAL_R_DURATION_CFG_ZQ_CAL_R_DURATION(32'h28)
        , .DDR_DDRC_CFG_ODT_POWERDOWN_CFG_ODT_POWERDOWN(32'h0), .DDR_DDRC_CFG_WL_CFG_WL(32'h8)
        , .DDR_DDRC_CFG_RL_CFG_RL(32'hE), .DDR_DDRC_CFG_BL_CFG_BL(32'h0)
        , .DDR_OPTIONS_TIP_CFG_PARAMS_ADDCMD_OFFSET(3'h7), .DDR_DDRC_CFG_ZQLATCH_DURATION_CFG_ZQLATCH_DURATION(32'h18)
        , .DDR_DDRC_CFG_ZQ_CAL_DURATION_CFG_ZQ_CAL_DURATION(32'h320), .DDR_DDRC_CFG_MRRI_CFG_MRRI(32'h12)
        , .DDR_DDRC_CFG_WR_POSTAMBLE_CFG_WR_POSTAMBLE(32'h0), .DDR_DDRC_CFG_SOC_ODT_CFG_SOC_ODT(32'h6)
        , .DDR_DDRC_CFG_ODTE_CK_CFG_ODTE_CK(32'h0), .DDR_DDRC_CFG_ODTE_CS_CFG_ODTE_CS(32'h0)
        , .DDR_DDRC_CFG_ODTD_CA_CFG_ODTD_CA(32'h0), .DDR_DDRC_CFG_RD_PREAMB_TOGGLE_CFG_RD_PREAMB_TOGGLE(32'h0)
        , .DDR_DDRC_CFG_RD_POSTAMBLE_CFG_RD_POSTAMBLE(32'h0), .DDR_DDRC_CFG_PU_CAL_CFG_PU_CAL(32'h0)
        , .DDR_DDRC_CFG_DQ_ODT_CFG_DQ_ODT(32'h2), .DDR_DDRC_CFG_CA_ODT_CFG_CA_ODT(32'h4)
        , .DDR_DDRC_CFG_MRD_CFG_MRD(32'hC), .DDR_DDRC_CFG_LPDDR4_FSP_OP_CFG_LPDDR4_FSP_OP(32'h1)
        , .CLK_MSS_SYS_CLOCK_CONFIG_CR_DIVIDER_CPU(2'h0), .CLK_MSS_SYS_CLOCK_CONFIG_CR_DIVIDER_AXI(2'h1)
        , .CLK_MSS_SYS_CLOCK_CONFIG_CR_DIVIDER_APB_AHB(2'h2), .CLK_MSS_CFM_PLL_CKMUX_PLL1_RFCLK0_SEL(2'h1)
        , .CLK_MSS_CFM_PLL_CKMUX_PLL1_RFCLK1_SEL(2'h1), .CLK_MSS_CFM_PLL_CKMUX_PLL0_RFCLK0_SEL(2'h1)
        , .CLK_MSS_CFM_PLL_CKMUX_PLL0_RFCLK1_SEL(2'h1), .CLK_MSS_CFM_PLL_CKMUX_CLK_IN_MAC_TSU_SEL(2'h1)
        , .SGMII_CLK_CNTL_REG_CLKMUX_PLL0_RFCLK0_SEL(2'h1), .SGMII_CLK_CNTL_REG_CLKMUX_PLL0_RFCLK1_SEL(2'h1)
        , .CLK_MSS_CFM_MSSCLKMUX_MSSCLK_MUX_SEL(2'h3), .CLK_MSS_CFM_MSSCLKMUX_CLK_STANDBY_SEL(1'h0)
        , .CLK_MSS_CFM_BCLKMUX_BCLK0_SEL(5'h8), .CLK_MSS_CFM_BCLKMUX_BCLK1_SEL(5'h10)
        , .CLK_MSS_CFM_BCLKMUX_BCLK2_SEL(5'h0), .CLK_MSS_CFM_BCLKMUX_BCLK3_SEL(5'h0)
        , .CLK_MSS_CFM_BCLKMUX_BCLK4_SEL(5'h0), .CLK_MSS_CFM_BCLKMUX_BCLK5_SEL(5'h0)
        , .CLK_MSS_PLL_PLL_CTRL_REG_RFCLK_SEL(1'h0), .CLK_SGMII_PLL_PLL_CTRL_REG_RFCLK_SEL(1'h0)
        , .CLK_DDR_PLL_PLL_CTRL_REG_RFCLK_SEL(1'h0), .DDR_MODEL_DDRPHY_MODE_DDRMODE(3'h4)
        , .DDR_MODEL_DDRPHY_MODE_POWER_DOWN(1'h0), .DDR_MODEL_DDRPHY_MODE_CRC(1'h0)
        , .DDR_MODEL_DDRPHY_MODE_ECC(1'h0), .DDR_MODEL_DDRPHY_MODE_BUS_WIDTH(3'h0)
        , .DDR_MODEL_DDRPHY_MODE_DMI_DBI(1'h0), .DDR_MODEL_DDRPHY_MODE_RANK(1'h0)
        , .DDR_MODEL_DDRPHY_MODE_DQ_DRIVE(2'h1), .DDR_MODEL_DDRPHY_MODE_DQS_DRIVE(2'h1)
        , .DDR_MODEL_DDRPHY_MODE_ADD_CMD_DRIVE(2'h2), .DDR_MODEL_DDRPHY_MODE_CLOCK_OUT_DRIVE(2'h2)
        , .DDR_IOBANK_RPC_ODT_DQ_RPC_ODT_DQ(32'h3), .DDR_IOBANK_RPC_ODT_DQS_RPC_ODT_DQS(32'h6)
        , .DDR_IOBANK_DPC_BITS_DPC_VRGEN_V(6'h10), .DDR_IOBANK_DPC_BITS_DPC_VRGEN_H(6'h2)
        , .DDR_IOBANK_DPC_BITS_DPC_VRGEN_EN_V(1'h1), .DDR_IOBANK_DPC_BITS_DPC_VRGEN_EN_H(1'h1)
        , .DDR_IOBANK_DPC_BITS_DPC_MOVE_EN_V(1'h0), .DDR_IOBANK_DPC_BITS_DPC_MOVE_EN_H(1'h0)
        , .DDR_IOBANK_DPC_BITS_DPC_VS(4'h2), .DDR_IOBANK_RPC_ODT_STATIC_DQ_RPC_ODT_STATIC_DQ(32'h5)
        , .DDR_IOBANK_RPC_ODT_STATIC_DQS_RPC_ODT_STATIC_DQS(32'h5), .DDR_IOBANK_RPC_ODT_STATIC_ADDCMD_RPC_ODT_STATIC_ADDCMD(32'h7)
        , .DDR_IOBANK_RPC_ODT_STATIC_CLKP_RPC_ODT_STATIC_CLKP(32'h7), .DDR_IOBANK_RPC_ODT_STATIC_CLKN_RPC_ODT_STATIC_CLKN(32'h7)
        , .DDR_IOBANK_RPC_IBUFMD_ADDCMD_RPC_IBUFMD_ADDCMD(32'h3), .DDR_IOBANK_RPC_IBUFMD_CLK_RPC_IBUFMD_CLK(32'h4)
        , .DDR_IOBANK_RPC_IBUFMD_DQ_RPC_IBUFMD_DQ(32'h3), .DDR_IOBANK_RPC_IBUFMD_DQS_RPC_IBUFMD_DQS(32'h4)
        , .DDR_IOBANK_RPC_SPARE0_DQ_RPC_SPARE0_DQ(32'h8000), .SGMII_SPARE_CNTL_REG_SPARE(32'hFF000000)
        , .TRACE_CR_ULTRASOC_FABRIC(1'b0), .MSS_IO_LOCKDOWN_CR_MSSIO_B2_LOCKDN_EN(1'b0)
        , .MSS_IO_LOCKDOWN_CR_MSSIO_B4_LOCKDN_EN(1'b0), .MSS_IO_LOCKDOWN_CR_SGMII_IO_LOCKDN_EN(1'b0)
        , .MSS_IO_LOCKDOWN_CR_DDR_IO_LOCKDN_EN(1'b0), .DLL0_CTRL0_PHASE_P(2'b11)
        , .DLL0_CTRL0_PHASE_S(2'b11), .DLL0_CTRL0_SEL_P(2'b00), .DLL0_CTRL0_SEL_S(2'b00)
        , .DLL0_CTRL0_REF_SEL(1'b0), .DLL0_CTRL0_FB_SEL(1'b0), .DLL0_CTRL0_DIV_SEL(1'b0)
        , .DLL0_CTRL0_ALU_UPD(2'b00), .DLL0_CTRL0_LOCK_FRC(1'b0), .DLL0_CTRL0_LOCK_FLT(2'b01)
        , .DLL0_CTRL0_LOCK_HIGH(4'b1000), .DLL0_CTRL0_LOCK_LOW(4'b1000)
        , .DLL0_CTRL1_SET_ALU(8'b00000000), .DLL0_CTRL1_ADJ_DEL4(7'b0000000)
        , .DLL0_CTRL1_TEST_S(1'b0), .DLL0_CTRL1_TEST_RING(1'b0), .DLL0_CTRL1_INIT_CODE(6'b000000)
        , .DLL0_CTRL1_RELOCK_FAST(1'b0), .DLL0_STAT0_RESET(1'b0), .DLL0_STAT0_BYPASS(1'b0)
        , .DLL0_STAT0_PHASE_MOVE_CLK(1'b1), .DLL1_CTRL0_PHASE_P(2'b11)
        , .DLL1_CTRL0_PHASE_S(2'b11), .DLL1_CTRL0_SEL_P(2'b00), .DLL1_CTRL0_SEL_S(2'b00)
        , .DLL1_CTRL0_REF_SEL(1'b0), .DLL1_CTRL0_FB_SEL(1'b0), .DLL1_CTRL0_DIV_SEL(1'b0)
        , .DLL1_CTRL0_ALU_UPD(2'b00), .DLL1_CTRL0_LOCK_FRC(1'b0), .DLL1_CTRL0_LOCK_FLT(2'b01)
        , .DLL1_CTRL0_LOCK_HIGH(4'b1000), .DLL1_CTRL0_LOCK_LOW(4'b1000)
        , .DLL1_CTRL1_SET_ALU(8'b00000000), .DLL1_CTRL1_ADJ_DEL4(7'b0000000)
        , .DLL1_CTRL1_TEST_S(1'b0), .DLL1_CTRL1_TEST_RING(1'b0), .DLL1_CTRL1_INIT_CODE(6'b000000)
        , .DLL1_CTRL1_RELOCK_FAST(1'b0), .DLL1_STAT0_RESET(1'b0), .DLL1_STAT0_BYPASS(1'b0)
        , .DLL1_STAT0_PHASE_MOVE_CLK(1'b1), .DLL2_CTRL0_PHASE_P(2'b11)
        , .DLL2_CTRL0_PHASE_S(2'b11), .DLL2_CTRL0_SEL_P(2'b00), .DLL2_CTRL0_SEL_S(2'b00)
        , .DLL2_CTRL0_REF_SEL(1'b0), .DLL2_CTRL0_FB_SEL(1'b0), .DLL2_CTRL0_DIV_SEL(1'b0)
        , .DLL2_CTRL0_ALU_UPD(2'b00), .DLL2_CTRL0_LOCK_FRC(1'b0), .DLL2_CTRL0_LOCK_FLT(2'b01)
        , .DLL2_CTRL0_LOCK_HIGH(4'b1000), .DLL2_CTRL0_LOCK_LOW(4'b1000)
        , .DLL2_CTRL1_SET_ALU(8'b00000000), .DLL2_CTRL1_ADJ_DEL4(7'b0000000)
        , .DLL2_CTRL1_TEST_S(1'b0), .DLL2_CTRL1_TEST_RING(1'b0), .DLL2_CTRL1_INIT_CODE(6'b000000)
        , .DLL2_CTRL1_RELOCK_FAST(1'b0), .DLL2_STAT0_RESET(1'b0), .DLL2_STAT0_BYPASS(1'b0)
        , .DLL2_STAT0_PHASE_MOVE_CLK(1'b1), .DLL3_CTRL0_PHASE_P(2'b11)
        , .DLL3_CTRL0_PHASE_S(2'b00), .DLL3_CTRL0_SEL_P(2'b00), .DLL3_CTRL0_SEL_S(2'b00)
        , .DLL3_CTRL0_REF_SEL(1'b0), .DLL3_CTRL0_FB_SEL(1'b0), .DLL3_CTRL0_DIV_SEL(1'b0)
        , .DLL3_CTRL0_ALU_UPD(2'b00), .DLL3_CTRL0_LOCK_FRC(1'b1), .DLL3_CTRL0_LOCK_FLT(2'b00)
        , .DLL3_CTRL0_LOCK_HIGH(4'b1000), .DLL3_CTRL0_LOCK_LOW(4'b1000)
        , .DLL3_CTRL1_SET_ALU(8'b10000000), .DLL3_CTRL1_ADJ_DEL4(7'b0000000)
        , .DLL3_CTRL1_TEST_S(1'b0), .DLL3_CTRL1_TEST_RING(1'b0), .DLL3_CTRL1_INIT_CODE(6'b000000)
        , .DLL3_CTRL1_RELOCK_FAST(1'b0), .DLL3_STAT0_RESET(1'b0), .DLL3_STAT0_BYPASS(1'b1)
        , .DLL3_STAT0_PHASE_MOVE_CLK(1'b1), .CRYPTO_SOFT_RESET_PERIPH(1'b1)
        , .CRYPTO_DLL_CTRL0_PHASE_P(2'b11), .CRYPTO_DLL_CTRL0_PHASE_S(2'b11)
        , .CRYPTO_DLL_CTRL0_SEL_P(2'b00), .CRYPTO_DLL_CTRL0_SEL_S(2'b00)
        , .CRYPTO_DLL_CTRL0_REF_SEL(1'b0), .CRYPTO_DLL_CTRL0_FB_SEL(1'b0)
        , .CRYPTO_DLL_CTRL0_DIV_SEL(1'b0), .CRYPTO_DLL_CTRL0_ALU_UPD(2'b00)
        , .CRYPTO_DLL_CTRL0_LOCK_FRC(1'b0), .CRYPTO_DLL_CTRL0_LOCK_FLT(2'b01)
        , .CRYPTO_DLL_CTRL0_LOCK_HIGH(4'b1000), .CRYPTO_DLL_CTRL0_LOCK_LOW(4'b1000)
        , .CRYPTO_DLL_CTRL1_SET_ALU(8'b00000000), .CRYPTO_DLL_CTRL1_ADJ_DEL4(7'b0000000)
        , .CRYPTO_DLL_CTRL1_TEST_S(1'b0), .CRYPTO_DLL_CTRL1_TEST_RING(1'b0)
        , .CRYPTO_DLL_CTRL1_INIT_CODE(6'b000000), .CRYPTO_DLL_CTRL1_RELOCK_FAST(1'b0)
        , .CRYPTO_DLL_STAT0_RESET(1'b0), .CRYPTO_DLL_STAT0_BYPASS(1'b0)
        , .CRYPTO_DLL_STAT0_PHASE_MOVE_CLK(1'b1), .CRYPTO_CONTROL_USER_SCB_CONTROL(1'b0)
        , .CRYPTO_CONTROL_USER_RESET(1'b0), .CRYPTO_CONTROL_USER_CLOCK_ENABLE(1'b1)
        , .CRYPTO_CONTROL_USER_CLOCK_SELECT(2'b01), .CRYPTO_CONTROL_USER_RAMS_ON(1'b1)
        , .CRYPTO_CONTROL_USER_DLL_ON(1'b1), .CRYPTO_CONTROL_USER_RING_OSC_ON(1'b1)
        , .CRYPTO_CONTROL_USER_PURGE(1'b0), .CRYPTO_CONTROL_USER_GO(1'b0)
        , .CRYPTO_INTERRUPT_ENABLE_COMPLETE(1'b0), .CRYPTO_INTERRUPT_ENABLE_ALARM(1'b0)
        , .CRYPTO_INTERRUPT_ENABLE_BUSERROR(1'b0), .CRYPTO_MARGIN_RAM(3'b000)
        , .CRYPTO_MARGIN_ROM(3'b000) )  I_MSS (.FIC_0_DLL_LOCK_M2F(
        FIC_0_DLL_LOCK_M2F), .FIC_1_DLL_LOCK_M2F(FIC_1_DLL_LOCK_M2F), 
        .FIC_2_DLL_LOCK_M2F(FIC_2_DLL_LOCK_M2F), .FIC_3_DLL_LOCK_M2F(
        FIC_3_DLL_LOCK_M2F), .FIC_0_AXI4_M_AWID({FIC_0_AXI4_M_AWID[7], 
        FIC_0_AXI4_M_AWID[6], FIC_0_AXI4_M_AWID[5], 
        FIC_0_AXI4_M_AWID[4], FIC_0_AXI4_M_AWID[3], 
        FIC_0_AXI4_M_AWID[2], FIC_0_AXI4_M_AWID[1], 
        FIC_0_AXI4_M_AWID[0]}), .FIC_0_AXI4_M_AWADDR({
        FIC_0_AXI4_M_AWADDR[37], FIC_0_AXI4_M_AWADDR[36], 
        FIC_0_AXI4_M_AWADDR[35], FIC_0_AXI4_M_AWADDR[34], 
        FIC_0_AXI4_M_AWADDR[33], FIC_0_AXI4_M_AWADDR[32], 
        FIC_0_AXI4_M_AWADDR[31], FIC_0_AXI4_M_AWADDR[30], 
        FIC_0_AXI4_M_AWADDR[29], FIC_0_AXI4_M_AWADDR[28], 
        FIC_0_AXI4_M_AWADDR[27], FIC_0_AXI4_M_AWADDR[26], 
        FIC_0_AXI4_M_AWADDR[25], FIC_0_AXI4_M_AWADDR[24], 
        FIC_0_AXI4_M_AWADDR[23], FIC_0_AXI4_M_AWADDR[22], 
        FIC_0_AXI4_M_AWADDR[21], FIC_0_AXI4_M_AWADDR[20], 
        FIC_0_AXI4_M_AWADDR[19], FIC_0_AXI4_M_AWADDR[18], 
        FIC_0_AXI4_M_AWADDR[17], FIC_0_AXI4_M_AWADDR[16], 
        FIC_0_AXI4_M_AWADDR[15], FIC_0_AXI4_M_AWADDR[14], 
        FIC_0_AXI4_M_AWADDR[13], FIC_0_AXI4_M_AWADDR[12], 
        FIC_0_AXI4_M_AWADDR[11], FIC_0_AXI4_M_AWADDR[10], 
        FIC_0_AXI4_M_AWADDR[9], FIC_0_AXI4_M_AWADDR[8], 
        FIC_0_AXI4_M_AWADDR[7], FIC_0_AXI4_M_AWADDR[6], 
        FIC_0_AXI4_M_AWADDR[5], FIC_0_AXI4_M_AWADDR[4], 
        FIC_0_AXI4_M_AWADDR[3], FIC_0_AXI4_M_AWADDR[2], 
        FIC_0_AXI4_M_AWADDR[1], FIC_0_AXI4_M_AWADDR[0]}), 
        .FIC_0_AXI4_M_AWLEN({FIC_0_AXI4_M_AWLEN[7], 
        FIC_0_AXI4_M_AWLEN[6], FIC_0_AXI4_M_AWLEN[5], 
        FIC_0_AXI4_M_AWLEN[4], FIC_0_AXI4_M_AWLEN[3], 
        FIC_0_AXI4_M_AWLEN[2], FIC_0_AXI4_M_AWLEN[1], 
        FIC_0_AXI4_M_AWLEN[0]}), .FIC_0_AXI4_M_AWSIZE({
        FIC_0_AXI4_M_AWSIZE[2], FIC_0_AXI4_M_AWSIZE[1], 
        FIC_0_AXI4_M_AWSIZE[0]}), .FIC_0_AXI4_M_AWBURST({
        FIC_0_AXI4_M_AWBURST[1], FIC_0_AXI4_M_AWBURST[0]}), 
        .FIC_0_AXI4_M_AWLOCK(FIC_0_AXI4_M_AWLOCK), .FIC_0_AXI4_M_AWQOS({
        FIC_0_AXI4_M_AWQOS[3], FIC_0_AXI4_M_AWQOS[2], 
        FIC_0_AXI4_M_AWQOS[1], FIC_0_AXI4_M_AWQOS[0]}), 
        .FIC_0_AXI4_M_AWCACHE({FIC_0_AXI4_M_AWCACHE[3], 
        FIC_0_AXI4_M_AWCACHE[2], FIC_0_AXI4_M_AWCACHE[1], 
        FIC_0_AXI4_M_AWCACHE[0]}), .FIC_0_AXI4_M_AWPROT({
        FIC_0_AXI4_M_AWPROT[2], FIC_0_AXI4_M_AWPROT[1], 
        FIC_0_AXI4_M_AWPROT[0]}), .FIC_0_AXI4_M_AWVALID(
        FIC_0_AXI4_M_AWVALID), .FIC_0_AXI4_M_WDATA({
        FIC_0_AXI4_M_WDATA[63], FIC_0_AXI4_M_WDATA[62], 
        FIC_0_AXI4_M_WDATA[61], FIC_0_AXI4_M_WDATA[60], 
        FIC_0_AXI4_M_WDATA[59], FIC_0_AXI4_M_WDATA[58], 
        FIC_0_AXI4_M_WDATA[57], FIC_0_AXI4_M_WDATA[56], 
        FIC_0_AXI4_M_WDATA[55], FIC_0_AXI4_M_WDATA[54], 
        FIC_0_AXI4_M_WDATA[53], FIC_0_AXI4_M_WDATA[52], 
        FIC_0_AXI4_M_WDATA[51], FIC_0_AXI4_M_WDATA[50], 
        FIC_0_AXI4_M_WDATA[49], FIC_0_AXI4_M_WDATA[48], 
        FIC_0_AXI4_M_WDATA[47], FIC_0_AXI4_M_WDATA[46], 
        FIC_0_AXI4_M_WDATA[45], FIC_0_AXI4_M_WDATA[44], 
        FIC_0_AXI4_M_WDATA[43], FIC_0_AXI4_M_WDATA[42], 
        FIC_0_AXI4_M_WDATA[41], FIC_0_AXI4_M_WDATA[40], 
        FIC_0_AXI4_M_WDATA[39], FIC_0_AXI4_M_WDATA[38], 
        FIC_0_AXI4_M_WDATA[37], FIC_0_AXI4_M_WDATA[36], 
        FIC_0_AXI4_M_WDATA[35], FIC_0_AXI4_M_WDATA[34], 
        FIC_0_AXI4_M_WDATA[33], FIC_0_AXI4_M_WDATA[32], 
        FIC_0_AXI4_M_WDATA[31], FIC_0_AXI4_M_WDATA[30], 
        FIC_0_AXI4_M_WDATA[29], FIC_0_AXI4_M_WDATA[28], 
        FIC_0_AXI4_M_WDATA[27], FIC_0_AXI4_M_WDATA[26], 
        FIC_0_AXI4_M_WDATA[25], FIC_0_AXI4_M_WDATA[24], 
        FIC_0_AXI4_M_WDATA[23], FIC_0_AXI4_M_WDATA[22], 
        FIC_0_AXI4_M_WDATA[21], FIC_0_AXI4_M_WDATA[20], 
        FIC_0_AXI4_M_WDATA[19], FIC_0_AXI4_M_WDATA[18], 
        FIC_0_AXI4_M_WDATA[17], FIC_0_AXI4_M_WDATA[16], 
        FIC_0_AXI4_M_WDATA[15], FIC_0_AXI4_M_WDATA[14], 
        FIC_0_AXI4_M_WDATA[13], FIC_0_AXI4_M_WDATA[12], 
        FIC_0_AXI4_M_WDATA[11], FIC_0_AXI4_M_WDATA[10], 
        FIC_0_AXI4_M_WDATA[9], FIC_0_AXI4_M_WDATA[8], 
        FIC_0_AXI4_M_WDATA[7], FIC_0_AXI4_M_WDATA[6], 
        FIC_0_AXI4_M_WDATA[5], FIC_0_AXI4_M_WDATA[4], 
        FIC_0_AXI4_M_WDATA[3], FIC_0_AXI4_M_WDATA[2], 
        FIC_0_AXI4_M_WDATA[1], FIC_0_AXI4_M_WDATA[0]}), 
        .FIC_0_AXI4_M_WSTRB({FIC_0_AXI4_M_WSTRB[7], 
        FIC_0_AXI4_M_WSTRB[6], FIC_0_AXI4_M_WSTRB[5], 
        FIC_0_AXI4_M_WSTRB[4], FIC_0_AXI4_M_WSTRB[3], 
        FIC_0_AXI4_M_WSTRB[2], FIC_0_AXI4_M_WSTRB[1], 
        FIC_0_AXI4_M_WSTRB[0]}), .FIC_0_AXI4_M_WLAST(
        FIC_0_AXI4_M_WLAST), .FIC_0_AXI4_M_WVALID(FIC_0_AXI4_M_WVALID), 
        .FIC_0_AXI4_M_BREADY(FIC_0_AXI4_M_BREADY), .FIC_0_AXI4_M_ARID({
        FIC_0_AXI4_M_ARID[7], FIC_0_AXI4_M_ARID[6], 
        FIC_0_AXI4_M_ARID[5], FIC_0_AXI4_M_ARID[4], 
        FIC_0_AXI4_M_ARID[3], FIC_0_AXI4_M_ARID[2], 
        FIC_0_AXI4_M_ARID[1], FIC_0_AXI4_M_ARID[0]}), 
        .FIC_0_AXI4_M_ARADDR({FIC_0_AXI4_M_ARADDR[37], 
        FIC_0_AXI4_M_ARADDR[36], FIC_0_AXI4_M_ARADDR[35], 
        FIC_0_AXI4_M_ARADDR[34], FIC_0_AXI4_M_ARADDR[33], 
        FIC_0_AXI4_M_ARADDR[32], FIC_0_AXI4_M_ARADDR[31], 
        FIC_0_AXI4_M_ARADDR[30], FIC_0_AXI4_M_ARADDR[29], 
        FIC_0_AXI4_M_ARADDR[28], FIC_0_AXI4_M_ARADDR[27], 
        FIC_0_AXI4_M_ARADDR[26], FIC_0_AXI4_M_ARADDR[25], 
        FIC_0_AXI4_M_ARADDR[24], FIC_0_AXI4_M_ARADDR[23], 
        FIC_0_AXI4_M_ARADDR[22], FIC_0_AXI4_M_ARADDR[21], 
        FIC_0_AXI4_M_ARADDR[20], FIC_0_AXI4_M_ARADDR[19], 
        FIC_0_AXI4_M_ARADDR[18], FIC_0_AXI4_M_ARADDR[17], 
        FIC_0_AXI4_M_ARADDR[16], FIC_0_AXI4_M_ARADDR[15], 
        FIC_0_AXI4_M_ARADDR[14], FIC_0_AXI4_M_ARADDR[13], 
        FIC_0_AXI4_M_ARADDR[12], FIC_0_AXI4_M_ARADDR[11], 
        FIC_0_AXI4_M_ARADDR[10], FIC_0_AXI4_M_ARADDR[9], 
        FIC_0_AXI4_M_ARADDR[8], FIC_0_AXI4_M_ARADDR[7], 
        FIC_0_AXI4_M_ARADDR[6], FIC_0_AXI4_M_ARADDR[5], 
        FIC_0_AXI4_M_ARADDR[4], FIC_0_AXI4_M_ARADDR[3], 
        FIC_0_AXI4_M_ARADDR[2], FIC_0_AXI4_M_ARADDR[1], 
        FIC_0_AXI4_M_ARADDR[0]}), .FIC_0_AXI4_M_ARLEN({
        FIC_0_AXI4_M_ARLEN[7], FIC_0_AXI4_M_ARLEN[6], 
        FIC_0_AXI4_M_ARLEN[5], FIC_0_AXI4_M_ARLEN[4], 
        FIC_0_AXI4_M_ARLEN[3], FIC_0_AXI4_M_ARLEN[2], 
        FIC_0_AXI4_M_ARLEN[1], FIC_0_AXI4_M_ARLEN[0]}), 
        .FIC_0_AXI4_M_ARSIZE({FIC_0_AXI4_M_ARSIZE[2], 
        FIC_0_AXI4_M_ARSIZE[1], FIC_0_AXI4_M_ARSIZE[0]}), 
        .FIC_0_AXI4_M_ARBURST({FIC_0_AXI4_M_ARBURST[1], 
        FIC_0_AXI4_M_ARBURST[0]}), .FIC_0_AXI4_M_ARLOCK(
        FIC_0_AXI4_M_ARLOCK), .FIC_0_AXI4_M_ARQOS({
        FIC_0_AXI4_M_ARQOS[3], FIC_0_AXI4_M_ARQOS[2], 
        FIC_0_AXI4_M_ARQOS[1], FIC_0_AXI4_M_ARQOS[0]}), 
        .FIC_0_AXI4_M_ARCACHE({FIC_0_AXI4_M_ARCACHE[3], 
        FIC_0_AXI4_M_ARCACHE[2], FIC_0_AXI4_M_ARCACHE[1], 
        FIC_0_AXI4_M_ARCACHE[0]}), .FIC_0_AXI4_M_ARPROT({
        FIC_0_AXI4_M_ARPROT[2], FIC_0_AXI4_M_ARPROT[1], 
        FIC_0_AXI4_M_ARPROT[0]}), .FIC_0_AXI4_M_ARVALID(
        FIC_0_AXI4_M_ARVALID), .FIC_0_AXI4_M_RREADY(
        FIC_0_AXI4_M_RREADY), .FIC_0_AXI4_S_AWREADY(
        FIC_0_AXI4_S_AWREADY), .FIC_0_AXI4_S_WREADY(
        FIC_0_AXI4_S_WREADY), .FIC_0_AXI4_S_BID({FIC_0_AXI4_S_BID[3], 
        FIC_0_AXI4_S_BID[2], FIC_0_AXI4_S_BID[1], FIC_0_AXI4_S_BID[0]})
        , .FIC_0_AXI4_S_BRESP({FIC_0_AXI4_S_BRESP[1], 
        FIC_0_AXI4_S_BRESP[0]}), .FIC_0_AXI4_S_BVALID(
        FIC_0_AXI4_S_BVALID), .FIC_0_AXI4_S_ARREADY(
        FIC_0_AXI4_S_ARREADY), .FIC_0_AXI4_S_RID({FIC_0_AXI4_S_RID[3], 
        FIC_0_AXI4_S_RID[2], FIC_0_AXI4_S_RID[1], FIC_0_AXI4_S_RID[0]})
        , .FIC_0_AXI4_S_RDATA({FIC_0_AXI4_S_RDATA[63], 
        FIC_0_AXI4_S_RDATA[62], FIC_0_AXI4_S_RDATA[61], 
        FIC_0_AXI4_S_RDATA[60], FIC_0_AXI4_S_RDATA[59], 
        FIC_0_AXI4_S_RDATA[58], FIC_0_AXI4_S_RDATA[57], 
        FIC_0_AXI4_S_RDATA[56], FIC_0_AXI4_S_RDATA[55], 
        FIC_0_AXI4_S_RDATA[54], FIC_0_AXI4_S_RDATA[53], 
        FIC_0_AXI4_S_RDATA[52], FIC_0_AXI4_S_RDATA[51], 
        FIC_0_AXI4_S_RDATA[50], FIC_0_AXI4_S_RDATA[49], 
        FIC_0_AXI4_S_RDATA[48], FIC_0_AXI4_S_RDATA[47], 
        FIC_0_AXI4_S_RDATA[46], FIC_0_AXI4_S_RDATA[45], 
        FIC_0_AXI4_S_RDATA[44], FIC_0_AXI4_S_RDATA[43], 
        FIC_0_AXI4_S_RDATA[42], FIC_0_AXI4_S_RDATA[41], 
        FIC_0_AXI4_S_RDATA[40], FIC_0_AXI4_S_RDATA[39], 
        FIC_0_AXI4_S_RDATA[38], FIC_0_AXI4_S_RDATA[37], 
        FIC_0_AXI4_S_RDATA[36], FIC_0_AXI4_S_RDATA[35], 
        FIC_0_AXI4_S_RDATA[34], FIC_0_AXI4_S_RDATA[33], 
        FIC_0_AXI4_S_RDATA[32], FIC_0_AXI4_S_RDATA[31], 
        FIC_0_AXI4_S_RDATA[30], FIC_0_AXI4_S_RDATA[29], 
        FIC_0_AXI4_S_RDATA[28], FIC_0_AXI4_S_RDATA[27], 
        FIC_0_AXI4_S_RDATA[26], FIC_0_AXI4_S_RDATA[25], 
        FIC_0_AXI4_S_RDATA[24], FIC_0_AXI4_S_RDATA[23], 
        FIC_0_AXI4_S_RDATA[22], FIC_0_AXI4_S_RDATA[21], 
        FIC_0_AXI4_S_RDATA[20], FIC_0_AXI4_S_RDATA[19], 
        FIC_0_AXI4_S_RDATA[18], FIC_0_AXI4_S_RDATA[17], 
        FIC_0_AXI4_S_RDATA[16], FIC_0_AXI4_S_RDATA[15], 
        FIC_0_AXI4_S_RDATA[14], FIC_0_AXI4_S_RDATA[13], 
        FIC_0_AXI4_S_RDATA[12], FIC_0_AXI4_S_RDATA[11], 
        FIC_0_AXI4_S_RDATA[10], FIC_0_AXI4_S_RDATA[9], 
        FIC_0_AXI4_S_RDATA[8], FIC_0_AXI4_S_RDATA[7], 
        FIC_0_AXI4_S_RDATA[6], FIC_0_AXI4_S_RDATA[5], 
        FIC_0_AXI4_S_RDATA[4], FIC_0_AXI4_S_RDATA[3], 
        FIC_0_AXI4_S_RDATA[2], FIC_0_AXI4_S_RDATA[1], 
        FIC_0_AXI4_S_RDATA[0]}), .FIC_0_AXI4_S_RRESP({
        FIC_0_AXI4_S_RRESP[1], FIC_0_AXI4_S_RRESP[0]}), 
        .FIC_0_AXI4_S_RLAST(FIC_0_AXI4_S_RLAST), .FIC_0_AXI4_S_RVALID(
        FIC_0_AXI4_S_RVALID), .FIC_1_AXI4_M_AWID({nc0, nc1, nc2, nc3, 
        nc4, nc5, nc6, nc7}), .FIC_1_AXI4_M_AWADDR({nc8, nc9, nc10, 
        nc11, nc12, nc13, nc14, nc15, nc16, nc17, nc18, nc19, nc20, 
        nc21, nc22, nc23, nc24, nc25, nc26, nc27, nc28, nc29, nc30, 
        nc31, nc32, nc33, nc34, nc35, nc36, nc37, nc38, nc39, nc40, 
        nc41, nc42, nc43, nc44, nc45}), .FIC_1_AXI4_M_AWLEN({nc46, 
        nc47, nc48, nc49, nc50, nc51, nc52, nc53}), 
        .FIC_1_AXI4_M_AWSIZE({nc54, nc55, nc56}), 
        .FIC_1_AXI4_M_AWBURST({nc57, nc58}), .FIC_1_AXI4_M_AWLOCK(), 
        .FIC_1_AXI4_M_AWQOS({nc59, nc60, nc61, nc62}), 
        .FIC_1_AXI4_M_AWCACHE({nc63, nc64, nc65, nc66}), 
        .FIC_1_AXI4_M_AWPROT({nc67, nc68, nc69}), 
        .FIC_1_AXI4_M_AWVALID(), .FIC_1_AXI4_M_WDATA({nc70, nc71, nc72, 
        nc73, nc74, nc75, nc76, nc77, nc78, nc79, nc80, nc81, nc82, 
        nc83, nc84, nc85, nc86, nc87, nc88, nc89, nc90, nc91, nc92, 
        nc93, nc94, nc95, nc96, nc97, nc98, nc99, nc100, nc101, nc102, 
        nc103, nc104, nc105, nc106, nc107, nc108, nc109, nc110, nc111, 
        nc112, nc113, nc114, nc115, nc116, nc117, nc118, nc119, nc120, 
        nc121, nc122, nc123, nc124, nc125, nc126, nc127, nc128, nc129, 
        nc130, nc131, nc132, nc133}), .FIC_1_AXI4_M_WSTRB({nc134, 
        nc135, nc136, nc137, nc138, nc139, nc140, nc141}), 
        .FIC_1_AXI4_M_WLAST(), .FIC_1_AXI4_M_WVALID(), 
        .FIC_1_AXI4_M_BREADY(), .FIC_1_AXI4_M_ARID({nc142, nc143, 
        nc144, nc145, nc146, nc147, nc148, nc149}), 
        .FIC_1_AXI4_M_ARADDR({nc150, nc151, nc152, nc153, nc154, nc155, 
        nc156, nc157, nc158, nc159, nc160, nc161, nc162, nc163, nc164, 
        nc165, nc166, nc167, nc168, nc169, nc170, nc171, nc172, nc173, 
        nc174, nc175, nc176, nc177, nc178, nc179, nc180, nc181, nc182, 
        nc183, nc184, nc185, nc186, nc187}), .FIC_1_AXI4_M_ARLEN({
        nc188, nc189, nc190, nc191, nc192, nc193, nc194, nc195}), 
        .FIC_1_AXI4_M_ARSIZE({nc196, nc197, nc198}), 
        .FIC_1_AXI4_M_ARBURST({nc199, nc200}), .FIC_1_AXI4_M_ARLOCK(), 
        .FIC_1_AXI4_M_ARQOS({nc201, nc202, nc203, nc204}), 
        .FIC_1_AXI4_M_ARCACHE({nc205, nc206, nc207, nc208}), 
        .FIC_1_AXI4_M_ARPROT({nc209, nc210, nc211}), 
        .FIC_1_AXI4_M_ARVALID(), .FIC_1_AXI4_M_RREADY(), 
        .FIC_1_AXI4_S_AWREADY(FIC_1_AXI4_S_AWREADY), 
        .FIC_1_AXI4_S_WREADY(FIC_1_AXI4_S_WREADY), .FIC_1_AXI4_S_BID({
        FIC_1_AXI4_S_BID[3], FIC_1_AXI4_S_BID[2], FIC_1_AXI4_S_BID[1], 
        FIC_1_AXI4_S_BID[0]}), .FIC_1_AXI4_S_BRESP({
        FIC_1_AXI4_S_BRESP[1], FIC_1_AXI4_S_BRESP[0]}), 
        .FIC_1_AXI4_S_BVALID(FIC_1_AXI4_S_BVALID), 
        .FIC_1_AXI4_S_ARREADY(FIC_1_AXI4_S_ARREADY), .FIC_1_AXI4_S_RID({
        FIC_1_AXI4_S_RID[3], FIC_1_AXI4_S_RID[2], FIC_1_AXI4_S_RID[1], 
        FIC_1_AXI4_S_RID[0]}), .FIC_1_AXI4_S_RDATA({
        FIC_1_AXI4_S_RDATA[63], FIC_1_AXI4_S_RDATA[62], 
        FIC_1_AXI4_S_RDATA[61], FIC_1_AXI4_S_RDATA[60], 
        FIC_1_AXI4_S_RDATA[59], FIC_1_AXI4_S_RDATA[58], 
        FIC_1_AXI4_S_RDATA[57], FIC_1_AXI4_S_RDATA[56], 
        FIC_1_AXI4_S_RDATA[55], FIC_1_AXI4_S_RDATA[54], 
        FIC_1_AXI4_S_RDATA[53], FIC_1_AXI4_S_RDATA[52], 
        FIC_1_AXI4_S_RDATA[51], FIC_1_AXI4_S_RDATA[50], 
        FIC_1_AXI4_S_RDATA[49], FIC_1_AXI4_S_RDATA[48], 
        FIC_1_AXI4_S_RDATA[47], FIC_1_AXI4_S_RDATA[46], 
        FIC_1_AXI4_S_RDATA[45], FIC_1_AXI4_S_RDATA[44], 
        FIC_1_AXI4_S_RDATA[43], FIC_1_AXI4_S_RDATA[42], 
        FIC_1_AXI4_S_RDATA[41], FIC_1_AXI4_S_RDATA[40], 
        FIC_1_AXI4_S_RDATA[39], FIC_1_AXI4_S_RDATA[38], 
        FIC_1_AXI4_S_RDATA[37], FIC_1_AXI4_S_RDATA[36], 
        FIC_1_AXI4_S_RDATA[35], FIC_1_AXI4_S_RDATA[34], 
        FIC_1_AXI4_S_RDATA[33], FIC_1_AXI4_S_RDATA[32], 
        FIC_1_AXI4_S_RDATA[31], FIC_1_AXI4_S_RDATA[30], 
        FIC_1_AXI4_S_RDATA[29], FIC_1_AXI4_S_RDATA[28], 
        FIC_1_AXI4_S_RDATA[27], FIC_1_AXI4_S_RDATA[26], 
        FIC_1_AXI4_S_RDATA[25], FIC_1_AXI4_S_RDATA[24], 
        FIC_1_AXI4_S_RDATA[23], FIC_1_AXI4_S_RDATA[22], 
        FIC_1_AXI4_S_RDATA[21], FIC_1_AXI4_S_RDATA[20], 
        FIC_1_AXI4_S_RDATA[19], FIC_1_AXI4_S_RDATA[18], 
        FIC_1_AXI4_S_RDATA[17], FIC_1_AXI4_S_RDATA[16], 
        FIC_1_AXI4_S_RDATA[15], FIC_1_AXI4_S_RDATA[14], 
        FIC_1_AXI4_S_RDATA[13], FIC_1_AXI4_S_RDATA[12], 
        FIC_1_AXI4_S_RDATA[11], FIC_1_AXI4_S_RDATA[10], 
        FIC_1_AXI4_S_RDATA[9], FIC_1_AXI4_S_RDATA[8], 
        FIC_1_AXI4_S_RDATA[7], FIC_1_AXI4_S_RDATA[6], 
        FIC_1_AXI4_S_RDATA[5], FIC_1_AXI4_S_RDATA[4], 
        FIC_1_AXI4_S_RDATA[3], FIC_1_AXI4_S_RDATA[2], 
        FIC_1_AXI4_S_RDATA[1], FIC_1_AXI4_S_RDATA[0]}), 
        .FIC_1_AXI4_S_RRESP({FIC_1_AXI4_S_RRESP[1], 
        FIC_1_AXI4_S_RRESP[0]}), .FIC_1_AXI4_S_RLAST(
        FIC_1_AXI4_S_RLAST), .FIC_1_AXI4_S_RVALID(FIC_1_AXI4_S_RVALID), 
        .FIC_2_AXI4_S_AWREADY(FIC_2_AXI4_S_AWREADY), 
        .FIC_2_AXI4_S_WREADY(FIC_2_AXI4_S_WREADY), .FIC_2_AXI4_S_BID({
        FIC_2_AXI4_S_BID[3], FIC_2_AXI4_S_BID[2], FIC_2_AXI4_S_BID[1], 
        FIC_2_AXI4_S_BID[0]}), .FIC_2_AXI4_S_BRESP({
        FIC_2_AXI4_S_BRESP[1], FIC_2_AXI4_S_BRESP[0]}), 
        .FIC_2_AXI4_S_BVALID(FIC_2_AXI4_S_BVALID), 
        .FIC_2_AXI4_S_ARREADY(FIC_2_AXI4_S_ARREADY), .FIC_2_AXI4_S_RID({
        FIC_2_AXI4_S_RID[3], FIC_2_AXI4_S_RID[2], FIC_2_AXI4_S_RID[1], 
        FIC_2_AXI4_S_RID[0]}), .FIC_2_AXI4_S_RDATA({
        FIC_2_AXI4_S_RDATA[63], FIC_2_AXI4_S_RDATA[62], 
        FIC_2_AXI4_S_RDATA[61], FIC_2_AXI4_S_RDATA[60], 
        FIC_2_AXI4_S_RDATA[59], FIC_2_AXI4_S_RDATA[58], 
        FIC_2_AXI4_S_RDATA[57], FIC_2_AXI4_S_RDATA[56], 
        FIC_2_AXI4_S_RDATA[55], FIC_2_AXI4_S_RDATA[54], 
        FIC_2_AXI4_S_RDATA[53], FIC_2_AXI4_S_RDATA[52], 
        FIC_2_AXI4_S_RDATA[51], FIC_2_AXI4_S_RDATA[50], 
        FIC_2_AXI4_S_RDATA[49], FIC_2_AXI4_S_RDATA[48], 
        FIC_2_AXI4_S_RDATA[47], FIC_2_AXI4_S_RDATA[46], 
        FIC_2_AXI4_S_RDATA[45], FIC_2_AXI4_S_RDATA[44], 
        FIC_2_AXI4_S_RDATA[43], FIC_2_AXI4_S_RDATA[42], 
        FIC_2_AXI4_S_RDATA[41], FIC_2_AXI4_S_RDATA[40], 
        FIC_2_AXI4_S_RDATA[39], FIC_2_AXI4_S_RDATA[38], 
        FIC_2_AXI4_S_RDATA[37], FIC_2_AXI4_S_RDATA[36], 
        FIC_2_AXI4_S_RDATA[35], FIC_2_AXI4_S_RDATA[34], 
        FIC_2_AXI4_S_RDATA[33], FIC_2_AXI4_S_RDATA[32], 
        FIC_2_AXI4_S_RDATA[31], FIC_2_AXI4_S_RDATA[30], 
        FIC_2_AXI4_S_RDATA[29], FIC_2_AXI4_S_RDATA[28], 
        FIC_2_AXI4_S_RDATA[27], FIC_2_AXI4_S_RDATA[26], 
        FIC_2_AXI4_S_RDATA[25], FIC_2_AXI4_S_RDATA[24], 
        FIC_2_AXI4_S_RDATA[23], FIC_2_AXI4_S_RDATA[22], 
        FIC_2_AXI4_S_RDATA[21], FIC_2_AXI4_S_RDATA[20], 
        FIC_2_AXI4_S_RDATA[19], FIC_2_AXI4_S_RDATA[18], 
        FIC_2_AXI4_S_RDATA[17], FIC_2_AXI4_S_RDATA[16], 
        FIC_2_AXI4_S_RDATA[15], FIC_2_AXI4_S_RDATA[14], 
        FIC_2_AXI4_S_RDATA[13], FIC_2_AXI4_S_RDATA[12], 
        FIC_2_AXI4_S_RDATA[11], FIC_2_AXI4_S_RDATA[10], 
        FIC_2_AXI4_S_RDATA[9], FIC_2_AXI4_S_RDATA[8], 
        FIC_2_AXI4_S_RDATA[7], FIC_2_AXI4_S_RDATA[6], 
        FIC_2_AXI4_S_RDATA[5], FIC_2_AXI4_S_RDATA[4], 
        FIC_2_AXI4_S_RDATA[3], FIC_2_AXI4_S_RDATA[2], 
        FIC_2_AXI4_S_RDATA[1], FIC_2_AXI4_S_RDATA[0]}), 
        .FIC_2_AXI4_S_RRESP({FIC_2_AXI4_S_RRESP[1], 
        FIC_2_AXI4_S_RRESP[0]}), .FIC_2_AXI4_S_RLAST(
        FIC_2_AXI4_S_RLAST), .FIC_2_AXI4_S_RVALID(FIC_2_AXI4_S_RVALID), 
        .FIC_3_APB_M_PSEL(FIC_3_APB_M_PSEL), .FIC_3_APB_M_PADDR({
        FIC_3_APB_M_PADDR[28], FIC_3_APB_M_PADDR[27], 
        FIC_3_APB_M_PADDR[26], FIC_3_APB_M_PADDR[25], 
        FIC_3_APB_M_PADDR[24], FIC_3_APB_M_PADDR[23], 
        FIC_3_APB_M_PADDR[22], FIC_3_APB_M_PADDR[21], 
        FIC_3_APB_M_PADDR[20], FIC_3_APB_M_PADDR[19], 
        FIC_3_APB_M_PADDR[18], FIC_3_APB_M_PADDR[17], 
        FIC_3_APB_M_PADDR[16], FIC_3_APB_M_PADDR[15], 
        FIC_3_APB_M_PADDR[14], FIC_3_APB_M_PADDR[13], 
        FIC_3_APB_M_PADDR[12], FIC_3_APB_M_PADDR[11], 
        FIC_3_APB_M_PADDR[10], FIC_3_APB_M_PADDR[9], 
        FIC_3_APB_M_PADDR[8], FIC_3_APB_M_PADDR[7], 
        FIC_3_APB_M_PADDR[6], FIC_3_APB_M_PADDR[5], 
        FIC_3_APB_M_PADDR[4], FIC_3_APB_M_PADDR[3], 
        FIC_3_APB_M_PADDR[2], FIC_3_APB_M_PADDR[1], 
        FIC_3_APB_M_PADDR[0]}), .FIC_3_APB_M_PWRITE(FIC_3_APB_M_PWRITE)
        , .FIC_3_APB_M_PENABLE(FIC_3_APB_M_PENABLE), 
        .FIC_3_APB_M_PSTRB({FIC_3_APB_M_PSTRB[3], FIC_3_APB_M_PSTRB[2], 
        FIC_3_APB_M_PSTRB[1], FIC_3_APB_M_PSTRB[0]}), 
        .FIC_3_APB_M_PWDATA({FIC_3_APB_M_PWDATA[31], 
        FIC_3_APB_M_PWDATA[30], FIC_3_APB_M_PWDATA[29], 
        FIC_3_APB_M_PWDATA[28], FIC_3_APB_M_PWDATA[27], 
        FIC_3_APB_M_PWDATA[26], FIC_3_APB_M_PWDATA[25], 
        FIC_3_APB_M_PWDATA[24], FIC_3_APB_M_PWDATA[23], 
        FIC_3_APB_M_PWDATA[22], FIC_3_APB_M_PWDATA[21], 
        FIC_3_APB_M_PWDATA[20], FIC_3_APB_M_PWDATA[19], 
        FIC_3_APB_M_PWDATA[18], FIC_3_APB_M_PWDATA[17], 
        FIC_3_APB_M_PWDATA[16], FIC_3_APB_M_PWDATA[15], 
        FIC_3_APB_M_PWDATA[14], FIC_3_APB_M_PWDATA[13], 
        FIC_3_APB_M_PWDATA[12], FIC_3_APB_M_PWDATA[11], 
        FIC_3_APB_M_PWDATA[10], FIC_3_APB_M_PWDATA[9], 
        FIC_3_APB_M_PWDATA[8], FIC_3_APB_M_PWDATA[7], 
        FIC_3_APB_M_PWDATA[6], FIC_3_APB_M_PWDATA[5], 
        FIC_3_APB_M_PWDATA[4], FIC_3_APB_M_PWDATA[3], 
        FIC_3_APB_M_PWDATA[2], FIC_3_APB_M_PWDATA[1], 
        FIC_3_APB_M_PWDATA[0]}), .MMUART_0_DTR_M2F(), 
        .MMUART_0_RTS_M2F(), .MMUART_0_TXD_M2F(MMUART_0_TXD_M2F), 
        .MMUART_0_TXD_OE_M2F(MMUART_0_TXD_OE_M2F), .MMUART_1_DTR_M2F(), 
        .MMUART_1_RTS_M2F(), .MMUART_1_TXD_M2F(MMUART_1_TXD_M2F), 
        .MMUART_1_TXD_OE_M2F(MMUART_1_TXD_OE_M2F), .MMUART_0_OUT1N_M2F(
        ), .MMUART_0_OUT2N_M2F(), .MMUART_0_TE_M2F(), 
        .MMUART_0_ESWM_M2F(), .MMUART_0_CLK_M2F(), 
        .MMUART_0_CLK_OE_M2F(), .MMUART_1_OUT1N_M2F(), 
        .MMUART_1_OUT2N_M2F(), .MMUART_1_TE_M2F(), .MMUART_1_ESWM_M2F()
        , .MMUART_1_CLK_M2F(), .MMUART_1_CLK_OE_M2F(), 
        .MMUART_2_TXD_M2F(MMUART_2_TXD_M2F), .MMUART_3_TXD_M2F(
        MMUART_3_TXD_M2F), .MMUART_4_TXD_M2F(MMUART_4_TXD_M2F), 
        .CAN_0_TX_EBL_M2F(CAN_0_TX_EBL_M2F), .CAN_0_TXBUS_M2F(
        CAN_0_TXBUS_M2F), .CAN_1_TX_EBL_M2F(), .CAN_1_TXBUS_M2F(), 
        .QSPI_SEL_M2F(), .QSPI_SEL_OE_M2F(), .QSPI_CLK_M2F(), 
        .QSPI_CLK_OE_M2F(), .QSPI_DATA_M2F({QSPI_DATA3_M2F, 
        QSPI_DATA2_M2F, nc212, nc213}), .QSPI_DATA_OE_M2F({
        QSPI_DATA3_OE_M2F, QSPI_DATA2_OE_M2F, nc214, nc215}), 
        .SPI_0_SS1_M2F(SPI_0_SS1_M2F), .SPI_0_SS1_OE_M2F(
        SPI_0_SS1_OE_M2F), .SPI_1_SS1_M2F(), .SPI_1_SS1_OE_M2F(), 
        .SPI_0_DO_M2F(SPI_0_DO_M2F), .SPI_0_DO_OE_M2F(SPI_0_DO_OE_M2F), 
        .SPI_0_CLK_M2F(SPI_0_CLK_M2F), .SPI_0_CLK_OE_M2F(
        SPI_0_CLK_OE_M2F), .SPI_1_DO_M2F(), .SPI_1_DO_OE_M2F(), 
        .SPI_1_CLK_M2F(), .SPI_1_CLK_OE_M2F(), .I2C_0_SCL_OE_M2F(
        I2C_0_SCL_OE_M2F_I_MSS_net), .I2C_0_SDA_OE_M2F(
        I2C_0_SDA_OE_M2F_I_MSS_net), .I2C_1_SCL_OE_M2F(), 
        .I2C_1_SDA_OE_M2F(), .I2C_0_SMBALERT_NO_M2F(), 
        .I2C_0_SMBSUS_NO_M2F(), .I2C_1_SMBALERT_NO_M2F(), 
        .I2C_1_SMBSUS_NO_M2F(), .GPIO_2_M2F({nc216, nc217, nc218, 
        GPIO_2_M2F_28, GPIO_2_M2F_27, GPIO_2_M2F_26, nc219, nc220, 
        nc221, nc222, nc223, nc224, GPIO_2_M2F_19, GPIO_2_M2F_18, 
        GPIO_2_M2F_17, GPIO_2_M2F_16, nc225, nc226, nc227, nc228, 
        nc229, nc230, nc231, nc232, nc233, nc234, nc235, nc236, nc237, 
        nc238, nc239, nc240}), .GPIO_2_OE_M2F({nc241, nc242, nc243, 
        nc244, nc245, nc246, nc247, nc248, nc249, nc250, nc251, nc252, 
        nc253, nc254, nc255, nc256, nc257, nc258, nc259, nc260, nc261, 
        nc262, nc263, nc264, nc265, nc266, nc267, nc268, nc269, nc270, 
        nc271, nc272}), .MAC_0_MDO_M2F(), .MAC_0_MDO_OE_M2F(), 
        .MAC_0_MDC_M2F(), .MAC_1_MDO_M2F(), .MAC_1_MDO_OE_M2F(), 
        .MAC_1_MDC_M2F(), .JTAG_TDO_M2F(), .JTAG_TDO_OE_M2F(), 
        .MSS_INT_M2F({MSS_INT_M2F[15], MSS_INT_M2F[14], 
        MSS_INT_M2F[13], MSS_INT_M2F[12], MSS_INT_M2F[11], 
        MSS_INT_M2F[10], MSS_INT_M2F[9], MSS_INT_M2F[8], 
        MSS_INT_M2F[7], MSS_INT_M2F[6], MSS_INT_M2F[5], MSS_INT_M2F[4], 
        MSS_INT_M2F[3], MSS_INT_M2F[2], MSS_INT_M2F[1], MSS_INT_M2F[0]})
        , .SPARE_M2F({nc273, nc274, nc275, nc276, nc277, nc278, nc279, 
        nc280, nc281, nc282, nc283, nc284, nc285, nc286, nc287, nc288, 
        nc289, nc290, nc291, nc292, nc293, nc294, nc295, nc296, nc297, 
        nc298, nc299, nc300, nc301, nc302, nc303, nc304, nc305, nc306, 
        nc307, nc308, nc309, nc310}), .PLL_CPU_LOCK_M2F(
        PLL_CPU_LOCK_M2F), .PLL_DDR_LOCK_M2F(PLL_DDR_LOCK_M2F), 
        .PLL_SGMII_LOCK_M2F(PLL_SGMII_LOCK_M2F), .MSS_STATUS_M2F({
        nc311, nc312, nc313, nc314, nc315, nc316, nc317, nc318, nc319, 
        nc320, nc321, nc322, nc323, nc324, nc325, nc326, nc327}), 
        .BOOT_FAIL_ERROR_M2F(), .MSS_RESET_N_M2F(MSS_RESET_N_M2F), 
        .SPARE_2_M2F({nc328, nc329, nc330, nc331, nc332}), 
        .SPARE_3_M2F(), .SPARE_4_M2F({nc333, nc334, nc335}), 
        .SPARE_5_M2F({nc336, nc337, nc338, nc339, nc340, nc341, nc342})
        , .WDOG_0_INTERRUPT_M2F(), .WDOG_1_INTERRUPT_M2F(), 
        .WDOG_2_INTERRUPT_M2F(), .WDOG_3_INTERRUPT_M2F(), 
        .WDOG_4_INTERRUPT_M2F(), .MPU_VIOLATION_FROM_FIC_0_M2F(), 
        .MPU_VIOLATION_FROM_FIC_1_M2F(), .MPU_VIOLATION_FROM_FIC_2_M2F(
        ), .MPU_VIOLATION_FROM_CRYPTO_M2F(), 
        .MPU_VIOLATION_FROM_MAC_0_M2F(), .MPU_VIOLATION_FROM_MAC_1_M2F(
        ), .MPU_VIOLATION_FROM_USB_M2F(), 
        .MPU_VIOLATION_FROM_EMMC_SD_M2F(), .MPU_VIOLATION_FROM_SCB_M2F(
        ), .MPU_VIOLATION_FROM_TRACE_M2F(), .REBOOT_REQUESTED_M2F(), 
        .CPU_IN_RESET_M2F(), .AXI_IN_RESET_M2F(), 
        .SCB_PERIPH_RESET_OCCURRED_M2F(), .SCB_MSS_RESET_OCCURRED_M2F()
        , .SCB_CPU_RESET_OCCURRED_M2F(), .DEBUGGER_RESET_OCCURRED_M2F()
        , .FABRIC_RESET_OCCURRED_M2F(), .WDOG_RESET_OCCURRED_M2F(), 
        .GPIO_RESET_OCCURRED_M2F(), .SCB_BUS_RESET_OCCURRED_M2F(), 
        .CPU_SOFT_RESET_OCCURRED_M2F(), .CPU_CLK_DIVIDER_M2F({nc343, 
        nc344}), .AXI_CLK_DIVIDER_M2F({nc345, nc346}), 
        .AHB_APB_CLK_DIVIDER_M2F({nc347, nc348}), 
        .USOC_CONTROL_DATA_M2F({nc349, nc350, nc351, nc352, nc353, 
        nc354, nc355, nc356}), .MAC_0_GMII_MII_TXD_M2F({nc357, nc358, 
        nc359, nc360, nc361, nc362, nc363, nc364}), 
        .MAC_0_GMII_MII_TX_EN_M2F(), .MAC_0_GMII_MII_TX_ER_M2F(), 
        .MAC_0_LOCAL_LOOPBACK_M2F(), .MAC_0_LOOPBACK_M2F(), 
        .MAC_0_HALF_DUPLEX_M2F(), .MAC_0_SPEED_MODE_M2F({nc365, nc366, 
        nc367, nc368}), .MAC_1_GMII_MII_TXD_M2F({nc369, nc370, nc371, 
        nc372, nc373, nc374, nc375, nc376}), .MAC_1_GMII_MII_TX_EN_M2F(
        ), .MAC_1_GMII_MII_TX_ER_M2F(), .MAC_1_LOCAL_LOOPBACK_M2F(), 
        .MAC_1_LOOPBACK_M2F(), .MAC_1_HALF_DUPLEX_M2F(), 
        .MAC_1_SPEED_MODE_M2F({nc377, nc378, nc379, nc380}), 
        .MAC_0_FILTER_DATA_M2F({nc381, nc382, nc383, nc384, nc385, 
        nc386, nc387, nc388, nc389, nc390, nc391, nc392, nc393, nc394, 
        nc395, nc396, nc397, nc398, nc399, nc400, nc401, nc402, nc403, 
        nc404, nc405, nc406, nc407, nc408, nc409, nc410, nc411, nc412, 
        nc413, nc414, nc415, nc416, nc417, nc418, nc419, nc420, nc421, 
        nc422, nc423, nc424, nc425, nc426, nc427, nc428, nc429, nc430, 
        nc431, nc432, nc433, nc434, nc435, nc436, nc437, nc438, nc439, 
        nc440, nc441, nc442, nc443, nc444, nc445, nc446, nc447, nc448, 
        nc449, nc450, nc451, nc452, nc453, nc454, nc455, nc456, nc457, 
        nc458, nc459, nc460, nc461, nc462, nc463, nc464, nc465, nc466, 
        nc467, nc468, nc469, nc470, nc471, nc472, nc473, nc474, nc475, 
        nc476, nc477, nc478, nc479, nc480, nc481, nc482, nc483, nc484, 
        nc485, nc486, nc487, nc488, nc489, nc490, nc491, nc492, nc493, 
        nc494, nc495, nc496, nc497, nc498, nc499, nc500, nc501, nc502, 
        nc503, nc504, nc505, nc506, nc507, nc508}), 
        .MAC_0_FILTER_SA_STB_M2F(), .MAC_0_FILTER_DA_STB_M2F(), 
        .MAC_0_FILTER_TYPE_STB_M2F(), .MAC_0_FILTER_VLAN_TAG1_STB_M2F()
        , .MAC_0_FILTER_VLAN_TAG2_STB_M2F(), 
        .MAC_0_FILTER_IP_SA_STB_M2F(), .MAC_0_FILTER_IP_DA_STB_M2F(), 
        .MAC_0_FILTER_SP_STB_M2F(), .MAC_0_FILTER_DP_STB_M2F(), 
        .MAC_0_FILTER_IPV6_M2F(), .MAC_0_WOL_M2F(), 
        .MAC_1_FILTER_DATA_M2F({nc509, nc510, nc511, nc512, nc513, 
        nc514, nc515, nc516, nc517, nc518, nc519, nc520, nc521, nc522, 
        nc523, nc524, nc525, nc526, nc527, nc528, nc529, nc530, nc531, 
        nc532, nc533, nc534, nc535, nc536, nc537, nc538, nc539, nc540, 
        nc541, nc542, nc543, nc544, nc545, nc546, nc547, nc548, nc549, 
        nc550, nc551, nc552, nc553, nc554, nc555, nc556, nc557, nc558, 
        nc559, nc560, nc561, nc562, nc563, nc564, nc565, nc566, nc567, 
        nc568, nc569, nc570, nc571, nc572, nc573, nc574, nc575, nc576, 
        nc577, nc578, nc579, nc580, nc581, nc582, nc583, nc584, nc585, 
        nc586, nc587, nc588, nc589, nc590, nc591, nc592, nc593, nc594, 
        nc595, nc596, nc597, nc598, nc599, nc600, nc601, nc602, nc603, 
        nc604, nc605, nc606, nc607, nc608, nc609, nc610, nc611, nc612, 
        nc613, nc614, nc615, nc616, nc617, nc618, nc619, nc620, nc621, 
        nc622, nc623, nc624, nc625, nc626, nc627, nc628, nc629, nc630, 
        nc631, nc632, nc633, nc634, nc635, nc636}), 
        .MAC_1_FILTER_SA_STB_M2F(), .MAC_1_FILTER_DA_STB_M2F(), 
        .MAC_1_FILTER_TYPE_STB_M2F(), .MAC_1_FILTER_VLAN_TAG1_STB_M2F()
        , .MAC_1_FILTER_VLAN_TAG2_STB_M2F(), 
        .MAC_1_FILTER_IP_SA_STB_M2F(), .MAC_1_FILTER_IP_DA_STB_M2F(), 
        .MAC_1_FILTER_SP_STB_M2F(), .MAC_1_FILTER_DP_STB_M2F(), 
        .MAC_1_FILTER_IPV6_M2F(), .MAC_1_WOL_M2F(), 
        .MAC_0_TSU_SOF_TX_M2F(MAC_0_TSU_SOF_TX_M2F), 
        .MAC_0_TSU_SYNC_FRAME_TX_M2F(MAC_0_TSU_SYNC_FRAME_TX_M2F), 
        .MAC_0_TSU_DELAY_REQ_TX_M2F(MAC_0_TSU_DELAY_REQ_TX_M2F), 
        .MAC_0_TSU_PDELAY_REQ_TX_M2F(MAC_0_TSU_PDELAY_REQ_TX_M2F), 
        .MAC_0_TSU_PDELAY_RESP_TX_M2F(MAC_0_TSU_PDELAY_RESP_TX_M2F), 
        .MAC_0_TSU_SOF_RX_M2F(MAC_0_TSU_SOF_RX_M2F), 
        .MAC_0_TSU_SYNC_FRAME_RX_M2F(MAC_0_TSU_SYNC_FRAME_RX_M2F), 
        .MAC_0_TSU_DELAY_REQ_RX_M2F(MAC_0_TSU_DELAY_REQ_RX_M2F), 
        .MAC_0_TSU_PDELAY_REQ_RX_M2F(MAC_0_TSU_PDELAY_REQ_RX_M2F), 
        .MAC_0_TSU_PDELAY_RESP_RX_M2F(MAC_0_TSU_PDELAY_RESP_RX_M2F), 
        .MAC_0_TSU_TIMER_CNT_M2F({MAC_0_TSU_TIMER_CNT_M2F[93], 
        MAC_0_TSU_TIMER_CNT_M2F[92], MAC_0_TSU_TIMER_CNT_M2F[91], 
        MAC_0_TSU_TIMER_CNT_M2F[90], MAC_0_TSU_TIMER_CNT_M2F[89], 
        MAC_0_TSU_TIMER_CNT_M2F[88], MAC_0_TSU_TIMER_CNT_M2F[87], 
        MAC_0_TSU_TIMER_CNT_M2F[86], MAC_0_TSU_TIMER_CNT_M2F[85], 
        MAC_0_TSU_TIMER_CNT_M2F[84], MAC_0_TSU_TIMER_CNT_M2F[83], 
        MAC_0_TSU_TIMER_CNT_M2F[82], MAC_0_TSU_TIMER_CNT_M2F[81], 
        MAC_0_TSU_TIMER_CNT_M2F[80], MAC_0_TSU_TIMER_CNT_M2F[79], 
        MAC_0_TSU_TIMER_CNT_M2F[78], MAC_0_TSU_TIMER_CNT_M2F[77], 
        MAC_0_TSU_TIMER_CNT_M2F[76], MAC_0_TSU_TIMER_CNT_M2F[75], 
        MAC_0_TSU_TIMER_CNT_M2F[74], MAC_0_TSU_TIMER_CNT_M2F[73], 
        MAC_0_TSU_TIMER_CNT_M2F[72], MAC_0_TSU_TIMER_CNT_M2F[71], 
        MAC_0_TSU_TIMER_CNT_M2F[70], MAC_0_TSU_TIMER_CNT_M2F[69], 
        MAC_0_TSU_TIMER_CNT_M2F[68], MAC_0_TSU_TIMER_CNT_M2F[67], 
        MAC_0_TSU_TIMER_CNT_M2F[66], MAC_0_TSU_TIMER_CNT_M2F[65], 
        MAC_0_TSU_TIMER_CNT_M2F[64], MAC_0_TSU_TIMER_CNT_M2F[63], 
        MAC_0_TSU_TIMER_CNT_M2F[62], MAC_0_TSU_TIMER_CNT_M2F[61], 
        MAC_0_TSU_TIMER_CNT_M2F[60], MAC_0_TSU_TIMER_CNT_M2F[59], 
        MAC_0_TSU_TIMER_CNT_M2F[58], MAC_0_TSU_TIMER_CNT_M2F[57], 
        MAC_0_TSU_TIMER_CNT_M2F[56], MAC_0_TSU_TIMER_CNT_M2F[55], 
        MAC_0_TSU_TIMER_CNT_M2F[54], MAC_0_TSU_TIMER_CNT_M2F[53], 
        MAC_0_TSU_TIMER_CNT_M2F[52], MAC_0_TSU_TIMER_CNT_M2F[51], 
        MAC_0_TSU_TIMER_CNT_M2F[50], MAC_0_TSU_TIMER_CNT_M2F[49], 
        MAC_0_TSU_TIMER_CNT_M2F[48], MAC_0_TSU_TIMER_CNT_M2F[47], 
        MAC_0_TSU_TIMER_CNT_M2F[46], MAC_0_TSU_TIMER_CNT_M2F[45], 
        MAC_0_TSU_TIMER_CNT_M2F[44], MAC_0_TSU_TIMER_CNT_M2F[43], 
        MAC_0_TSU_TIMER_CNT_M2F[42], MAC_0_TSU_TIMER_CNT_M2F[41], 
        MAC_0_TSU_TIMER_CNT_M2F[40], MAC_0_TSU_TIMER_CNT_M2F[39], 
        MAC_0_TSU_TIMER_CNT_M2F[38], MAC_0_TSU_TIMER_CNT_M2F[37], 
        MAC_0_TSU_TIMER_CNT_M2F[36], MAC_0_TSU_TIMER_CNT_M2F[35], 
        MAC_0_TSU_TIMER_CNT_M2F[34], MAC_0_TSU_TIMER_CNT_M2F[33], 
        MAC_0_TSU_TIMER_CNT_M2F[32], MAC_0_TSU_TIMER_CNT_M2F[31], 
        MAC_0_TSU_TIMER_CNT_M2F[30], MAC_0_TSU_TIMER_CNT_M2F[29], 
        MAC_0_TSU_TIMER_CNT_M2F[28], MAC_0_TSU_TIMER_CNT_M2F[27], 
        MAC_0_TSU_TIMER_CNT_M2F[26], MAC_0_TSU_TIMER_CNT_M2F[25], 
        MAC_0_TSU_TIMER_CNT_M2F[24], MAC_0_TSU_TIMER_CNT_M2F[23], 
        MAC_0_TSU_TIMER_CNT_M2F[22], MAC_0_TSU_TIMER_CNT_M2F[21], 
        MAC_0_TSU_TIMER_CNT_M2F[20], MAC_0_TSU_TIMER_CNT_M2F[19], 
        MAC_0_TSU_TIMER_CNT_M2F[18], MAC_0_TSU_TIMER_CNT_M2F[17], 
        MAC_0_TSU_TIMER_CNT_M2F[16], MAC_0_TSU_TIMER_CNT_M2F[15], 
        MAC_0_TSU_TIMER_CNT_M2F[14], MAC_0_TSU_TIMER_CNT_M2F[13], 
        MAC_0_TSU_TIMER_CNT_M2F[12], MAC_0_TSU_TIMER_CNT_M2F[11], 
        MAC_0_TSU_TIMER_CNT_M2F[10], MAC_0_TSU_TIMER_CNT_M2F[9], 
        MAC_0_TSU_TIMER_CNT_M2F[8], MAC_0_TSU_TIMER_CNT_M2F[7], 
        MAC_0_TSU_TIMER_CNT_M2F[6], MAC_0_TSU_TIMER_CNT_M2F[5], 
        MAC_0_TSU_TIMER_CNT_M2F[4], MAC_0_TSU_TIMER_CNT_M2F[3], 
        MAC_0_TSU_TIMER_CNT_M2F[2], MAC_0_TSU_TIMER_CNT_M2F[1], 
        MAC_0_TSU_TIMER_CNT_M2F[0]}), .MAC_0_TSU_TIMER_CMP_VAL_M2F(), 
        .MAC_1_TSU_SOF_TX_M2F(MAC_1_TSU_SOF_TX_M2F), 
        .MAC_1_TSU_SYNC_FRAME_TX_M2F(MAC_1_TSU_SYNC_FRAME_TX_M2F), 
        .MAC_1_TSU_DELAY_REQ_TX_M2F(MAC_1_TSU_DELAY_REQ_TX_M2F), 
        .MAC_1_TSU_PDELAY_REQ_TX_M2F(MAC_1_TSU_PDELAY_REQ_TX_M2F), 
        .MAC_1_TSU_PDELAY_RESP_TX_M2F(MAC_1_TSU_PDELAY_RESP_TX_M2F), 
        .MAC_1_TSU_SOF_RX_M2F(MAC_1_TSU_SOF_RX_M2F), 
        .MAC_1_TSU_SYNC_FRAME_RX_M2F(MAC_1_TSU_SYNC_FRAME_RX_M2F), 
        .MAC_1_TSU_DELAY_REQ_RX_M2F(MAC_1_TSU_DELAY_REQ_RX_M2F), 
        .MAC_1_TSU_PDELAY_REQ_RX_M2F(MAC_1_TSU_PDELAY_REQ_RX_M2F), 
        .MAC_1_TSU_PDELAY_RESP_RX_M2F(MAC_1_TSU_PDELAY_RESP_RX_M2F), 
        .MAC_1_TSU_TIMER_CNT_M2F({MAC_1_TSU_TIMER_CNT_M2F[93], 
        MAC_1_TSU_TIMER_CNT_M2F[92], MAC_1_TSU_TIMER_CNT_M2F[91], 
        MAC_1_TSU_TIMER_CNT_M2F[90], MAC_1_TSU_TIMER_CNT_M2F[89], 
        MAC_1_TSU_TIMER_CNT_M2F[88], MAC_1_TSU_TIMER_CNT_M2F[87], 
        MAC_1_TSU_TIMER_CNT_M2F[86], MAC_1_TSU_TIMER_CNT_M2F[85], 
        MAC_1_TSU_TIMER_CNT_M2F[84], MAC_1_TSU_TIMER_CNT_M2F[83], 
        MAC_1_TSU_TIMER_CNT_M2F[82], MAC_1_TSU_TIMER_CNT_M2F[81], 
        MAC_1_TSU_TIMER_CNT_M2F[80], MAC_1_TSU_TIMER_CNT_M2F[79], 
        MAC_1_TSU_TIMER_CNT_M2F[78], MAC_1_TSU_TIMER_CNT_M2F[77], 
        MAC_1_TSU_TIMER_CNT_M2F[76], MAC_1_TSU_TIMER_CNT_M2F[75], 
        MAC_1_TSU_TIMER_CNT_M2F[74], MAC_1_TSU_TIMER_CNT_M2F[73], 
        MAC_1_TSU_TIMER_CNT_M2F[72], MAC_1_TSU_TIMER_CNT_M2F[71], 
        MAC_1_TSU_TIMER_CNT_M2F[70], MAC_1_TSU_TIMER_CNT_M2F[69], 
        MAC_1_TSU_TIMER_CNT_M2F[68], MAC_1_TSU_TIMER_CNT_M2F[67], 
        MAC_1_TSU_TIMER_CNT_M2F[66], MAC_1_TSU_TIMER_CNT_M2F[65], 
        MAC_1_TSU_TIMER_CNT_M2F[64], MAC_1_TSU_TIMER_CNT_M2F[63], 
        MAC_1_TSU_TIMER_CNT_M2F[62], MAC_1_TSU_TIMER_CNT_M2F[61], 
        MAC_1_TSU_TIMER_CNT_M2F[60], MAC_1_TSU_TIMER_CNT_M2F[59], 
        MAC_1_TSU_TIMER_CNT_M2F[58], MAC_1_TSU_TIMER_CNT_M2F[57], 
        MAC_1_TSU_TIMER_CNT_M2F[56], MAC_1_TSU_TIMER_CNT_M2F[55], 
        MAC_1_TSU_TIMER_CNT_M2F[54], MAC_1_TSU_TIMER_CNT_M2F[53], 
        MAC_1_TSU_TIMER_CNT_M2F[52], MAC_1_TSU_TIMER_CNT_M2F[51], 
        MAC_1_TSU_TIMER_CNT_M2F[50], MAC_1_TSU_TIMER_CNT_M2F[49], 
        MAC_1_TSU_TIMER_CNT_M2F[48], MAC_1_TSU_TIMER_CNT_M2F[47], 
        MAC_1_TSU_TIMER_CNT_M2F[46], MAC_1_TSU_TIMER_CNT_M2F[45], 
        MAC_1_TSU_TIMER_CNT_M2F[44], MAC_1_TSU_TIMER_CNT_M2F[43], 
        MAC_1_TSU_TIMER_CNT_M2F[42], MAC_1_TSU_TIMER_CNT_M2F[41], 
        MAC_1_TSU_TIMER_CNT_M2F[40], MAC_1_TSU_TIMER_CNT_M2F[39], 
        MAC_1_TSU_TIMER_CNT_M2F[38], MAC_1_TSU_TIMER_CNT_M2F[37], 
        MAC_1_TSU_TIMER_CNT_M2F[36], MAC_1_TSU_TIMER_CNT_M2F[35], 
        MAC_1_TSU_TIMER_CNT_M2F[34], MAC_1_TSU_TIMER_CNT_M2F[33], 
        MAC_1_TSU_TIMER_CNT_M2F[32], MAC_1_TSU_TIMER_CNT_M2F[31], 
        MAC_1_TSU_TIMER_CNT_M2F[30], MAC_1_TSU_TIMER_CNT_M2F[29], 
        MAC_1_TSU_TIMER_CNT_M2F[28], MAC_1_TSU_TIMER_CNT_M2F[27], 
        MAC_1_TSU_TIMER_CNT_M2F[26], MAC_1_TSU_TIMER_CNT_M2F[25], 
        MAC_1_TSU_TIMER_CNT_M2F[24], MAC_1_TSU_TIMER_CNT_M2F[23], 
        MAC_1_TSU_TIMER_CNT_M2F[22], MAC_1_TSU_TIMER_CNT_M2F[21], 
        MAC_1_TSU_TIMER_CNT_M2F[20], MAC_1_TSU_TIMER_CNT_M2F[19], 
        MAC_1_TSU_TIMER_CNT_M2F[18], MAC_1_TSU_TIMER_CNT_M2F[17], 
        MAC_1_TSU_TIMER_CNT_M2F[16], MAC_1_TSU_TIMER_CNT_M2F[15], 
        MAC_1_TSU_TIMER_CNT_M2F[14], MAC_1_TSU_TIMER_CNT_M2F[13], 
        MAC_1_TSU_TIMER_CNT_M2F[12], MAC_1_TSU_TIMER_CNT_M2F[11], 
        MAC_1_TSU_TIMER_CNT_M2F[10], MAC_1_TSU_TIMER_CNT_M2F[9], 
        MAC_1_TSU_TIMER_CNT_M2F[8], MAC_1_TSU_TIMER_CNT_M2F[7], 
        MAC_1_TSU_TIMER_CNT_M2F[6], MAC_1_TSU_TIMER_CNT_M2F[5], 
        MAC_1_TSU_TIMER_CNT_M2F[4], MAC_1_TSU_TIMER_CNT_M2F[3], 
        MAC_1_TSU_TIMER_CNT_M2F[2], MAC_1_TSU_TIMER_CNT_M2F[1], 
        MAC_1_TSU_TIMER_CNT_M2F[0]}), .MAC_1_TSU_TIMER_CMP_VAL_M2F(), 
        .CRYPTO_DLL_LOCK_M2F(), .CRYPTO_AHB_M_HADDR({nc637, nc638, 
        nc639, nc640, nc641, nc642, nc643, nc644, nc645, nc646, nc647, 
        nc648, nc649, nc650, nc651, nc652, nc653, nc654, nc655, nc656, 
        nc657, nc658, nc659, nc660, nc661, nc662, nc663, nc664, nc665, 
        nc666, nc667, nc668}), .CRYPTO_AHB_M_HWDATA({nc669, nc670, 
        nc671, nc672, nc673, nc674, nc675, nc676, nc677, nc678, nc679, 
        nc680, nc681, nc682, nc683, nc684, nc685, nc686, nc687, nc688, 
        nc689, nc690, nc691, nc692, nc693, nc694, nc695, nc696, nc697, 
        nc698, nc699, nc700}), .CRYPTO_AHB_M_HSIZE({nc701, nc702}), 
        .CRYPTO_AHB_M_HTRANS({nc703, nc704}), .CRYPTO_AHB_M_HWRITE(), 
        .CRYPTO_AHB_M_HMASTLOCK(), .CRYPTO_AHB_S_HREADYOUT(), 
        .CRYPTO_AHB_S_HRESP(), .CRYPTO_AHB_S_HRDATA({nc705, nc706, 
        nc707, nc708, nc709, nc710, nc711, nc712, nc713, nc714, nc715, 
        nc716, nc717, nc718, nc719, nc720, nc721, nc722, nc723, nc724, 
        nc725, nc726, nc727, nc728, nc729, nc730, nc731, nc732, nc733, 
        nc734, nc735, nc736}), .CRYPTO_BUSY_M2F(), 
        .CRYPTO_COMPLETE_M2F(), .CRYPTO_ALARM_M2F(), 
        .CRYPTO_BUSERROR_M2F(), .CRYPTO_MSS_REQUEST_M2F(), 
        .CRYPTO_MSS_RELEASE_M2F(), .CRYPTO_OWNER_M2F(), 
        .CRYPTO_MSS_OWNER_M2F(), .CRYPTO_XWADDR_M2F({nc737, nc738, 
        nc739, nc740, nc741, nc742, nc743, nc744, nc745, nc746}), 
        .CRYPTO_XINACCEPT_M2F(), .CRYPTO_XRDATA_M2F({nc747, nc748, 
        nc749, nc750, nc751, nc752, nc753, nc754, nc755, nc756, nc757, 
        nc758, nc759, nc760, nc761, nc762, nc763, nc764, nc765, nc766, 
        nc767, nc768, nc769, nc770, nc771, nc772, nc773, nc774, nc775, 
        nc776, nc777, nc778}), .CRYPTO_XRADDR_M2F({nc779, nc780, nc781, 
        nc782, nc783, nc784, nc785, nc786, nc787, nc788}), 
        .CRYPTO_XVALIDOUT_M2F(), .CRYPTO_MESH_ERROR_M2F(), .FIC_0_ACLK(
        FIC_0_ACLK), .FIC_0_AXI4_M_AWREADY(FIC_0_AXI4_M_AWREADY), 
        .FIC_0_AXI4_M_WREADY(FIC_0_AXI4_M_WREADY), .FIC_0_AXI4_M_BID({
        FIC_0_AXI4_M_BID[7], FIC_0_AXI4_M_BID[6], FIC_0_AXI4_M_BID[5], 
        FIC_0_AXI4_M_BID[4], FIC_0_AXI4_M_BID[3], FIC_0_AXI4_M_BID[2], 
        FIC_0_AXI4_M_BID[1], FIC_0_AXI4_M_BID[0]}), 
        .FIC_0_AXI4_M_BRESP({FIC_0_AXI4_M_BRESP[1], 
        FIC_0_AXI4_M_BRESP[0]}), .FIC_0_AXI4_M_BVALID(
        FIC_0_AXI4_M_BVALID), .FIC_0_AXI4_M_ARREADY(
        FIC_0_AXI4_M_ARREADY), .FIC_0_AXI4_M_RID({FIC_0_AXI4_M_RID[7], 
        FIC_0_AXI4_M_RID[6], FIC_0_AXI4_M_RID[5], FIC_0_AXI4_M_RID[4], 
        FIC_0_AXI4_M_RID[3], FIC_0_AXI4_M_RID[2], FIC_0_AXI4_M_RID[1], 
        FIC_0_AXI4_M_RID[0]}), .FIC_0_AXI4_M_RDATA({
        FIC_0_AXI4_M_RDATA[63], FIC_0_AXI4_M_RDATA[62], 
        FIC_0_AXI4_M_RDATA[61], FIC_0_AXI4_M_RDATA[60], 
        FIC_0_AXI4_M_RDATA[59], FIC_0_AXI4_M_RDATA[58], 
        FIC_0_AXI4_M_RDATA[57], FIC_0_AXI4_M_RDATA[56], 
        FIC_0_AXI4_M_RDATA[55], FIC_0_AXI4_M_RDATA[54], 
        FIC_0_AXI4_M_RDATA[53], FIC_0_AXI4_M_RDATA[52], 
        FIC_0_AXI4_M_RDATA[51], FIC_0_AXI4_M_RDATA[50], 
        FIC_0_AXI4_M_RDATA[49], FIC_0_AXI4_M_RDATA[48], 
        FIC_0_AXI4_M_RDATA[47], FIC_0_AXI4_M_RDATA[46], 
        FIC_0_AXI4_M_RDATA[45], FIC_0_AXI4_M_RDATA[44], 
        FIC_0_AXI4_M_RDATA[43], FIC_0_AXI4_M_RDATA[42], 
        FIC_0_AXI4_M_RDATA[41], FIC_0_AXI4_M_RDATA[40], 
        FIC_0_AXI4_M_RDATA[39], FIC_0_AXI4_M_RDATA[38], 
        FIC_0_AXI4_M_RDATA[37], FIC_0_AXI4_M_RDATA[36], 
        FIC_0_AXI4_M_RDATA[35], FIC_0_AXI4_M_RDATA[34], 
        FIC_0_AXI4_M_RDATA[33], FIC_0_AXI4_M_RDATA[32], 
        FIC_0_AXI4_M_RDATA[31], FIC_0_AXI4_M_RDATA[30], 
        FIC_0_AXI4_M_RDATA[29], FIC_0_AXI4_M_RDATA[28], 
        FIC_0_AXI4_M_RDATA[27], FIC_0_AXI4_M_RDATA[26], 
        FIC_0_AXI4_M_RDATA[25], FIC_0_AXI4_M_RDATA[24], 
        FIC_0_AXI4_M_RDATA[23], FIC_0_AXI4_M_RDATA[22], 
        FIC_0_AXI4_M_RDATA[21], FIC_0_AXI4_M_RDATA[20], 
        FIC_0_AXI4_M_RDATA[19], FIC_0_AXI4_M_RDATA[18], 
        FIC_0_AXI4_M_RDATA[17], FIC_0_AXI4_M_RDATA[16], 
        FIC_0_AXI4_M_RDATA[15], FIC_0_AXI4_M_RDATA[14], 
        FIC_0_AXI4_M_RDATA[13], FIC_0_AXI4_M_RDATA[12], 
        FIC_0_AXI4_M_RDATA[11], FIC_0_AXI4_M_RDATA[10], 
        FIC_0_AXI4_M_RDATA[9], FIC_0_AXI4_M_RDATA[8], 
        FIC_0_AXI4_M_RDATA[7], FIC_0_AXI4_M_RDATA[6], 
        FIC_0_AXI4_M_RDATA[5], FIC_0_AXI4_M_RDATA[4], 
        FIC_0_AXI4_M_RDATA[3], FIC_0_AXI4_M_RDATA[2], 
        FIC_0_AXI4_M_RDATA[1], FIC_0_AXI4_M_RDATA[0]}), 
        .FIC_0_AXI4_M_RRESP({FIC_0_AXI4_M_RRESP[1], 
        FIC_0_AXI4_M_RRESP[0]}), .FIC_0_AXI4_M_RLAST(
        FIC_0_AXI4_M_RLAST), .FIC_0_AXI4_M_RVALID(FIC_0_AXI4_M_RVALID), 
        .FIC_0_AXI4_S_AWID({FIC_0_AXI4_S_AWID[3], FIC_0_AXI4_S_AWID[2], 
        FIC_0_AXI4_S_AWID[1], FIC_0_AXI4_S_AWID[0]}), 
        .FIC_0_AXI4_S_AWADDR({FIC_0_AXI4_S_AWADDR[37], 
        FIC_0_AXI4_S_AWADDR[36], FIC_0_AXI4_S_AWADDR[35], 
        FIC_0_AXI4_S_AWADDR[34], FIC_0_AXI4_S_AWADDR[33], 
        FIC_0_AXI4_S_AWADDR[32], FIC_0_AXI4_S_AWADDR[31], 
        FIC_0_AXI4_S_AWADDR[30], FIC_0_AXI4_S_AWADDR[29], 
        FIC_0_AXI4_S_AWADDR[28], FIC_0_AXI4_S_AWADDR[27], 
        FIC_0_AXI4_S_AWADDR[26], FIC_0_AXI4_S_AWADDR[25], 
        FIC_0_AXI4_S_AWADDR[24], FIC_0_AXI4_S_AWADDR[23], 
        FIC_0_AXI4_S_AWADDR[22], FIC_0_AXI4_S_AWADDR[21], 
        FIC_0_AXI4_S_AWADDR[20], FIC_0_AXI4_S_AWADDR[19], 
        FIC_0_AXI4_S_AWADDR[18], FIC_0_AXI4_S_AWADDR[17], 
        FIC_0_AXI4_S_AWADDR[16], FIC_0_AXI4_S_AWADDR[15], 
        FIC_0_AXI4_S_AWADDR[14], FIC_0_AXI4_S_AWADDR[13], 
        FIC_0_AXI4_S_AWADDR[12], FIC_0_AXI4_S_AWADDR[11], 
        FIC_0_AXI4_S_AWADDR[10], FIC_0_AXI4_S_AWADDR[9], 
        FIC_0_AXI4_S_AWADDR[8], FIC_0_AXI4_S_AWADDR[7], 
        FIC_0_AXI4_S_AWADDR[6], FIC_0_AXI4_S_AWADDR[5], 
        FIC_0_AXI4_S_AWADDR[4], FIC_0_AXI4_S_AWADDR[3], 
        FIC_0_AXI4_S_AWADDR[2], FIC_0_AXI4_S_AWADDR[1], 
        FIC_0_AXI4_S_AWADDR[0]}), .FIC_0_AXI4_S_AWLEN({
        FIC_0_AXI4_S_AWLEN[7], FIC_0_AXI4_S_AWLEN[6], 
        FIC_0_AXI4_S_AWLEN[5], FIC_0_AXI4_S_AWLEN[4], 
        FIC_0_AXI4_S_AWLEN[3], FIC_0_AXI4_S_AWLEN[2], 
        FIC_0_AXI4_S_AWLEN[1], FIC_0_AXI4_S_AWLEN[0]}), 
        .FIC_0_AXI4_S_AWSIZE({FIC_0_AXI4_S_AWSIZE[2], 
        FIC_0_AXI4_S_AWSIZE[1], FIC_0_AXI4_S_AWSIZE[0]}), 
        .FIC_0_AXI4_S_AWBURST({FIC_0_AXI4_S_AWBURST[1], 
        FIC_0_AXI4_S_AWBURST[0]}), .FIC_0_AXI4_S_AWQOS({
        FIC_0_AXI4_S_AWQOS[3], FIC_0_AXI4_S_AWQOS[2], 
        FIC_0_AXI4_S_AWQOS[1], FIC_0_AXI4_S_AWQOS[0]}), 
        .FIC_0_AXI4_S_AWLOCK(FIC_0_AXI4_S_AWLOCK), 
        .FIC_0_AXI4_S_AWCACHE({FIC_0_AXI4_S_AWCACHE[3], 
        FIC_0_AXI4_S_AWCACHE[2], FIC_0_AXI4_S_AWCACHE[1], 
        FIC_0_AXI4_S_AWCACHE[0]}), .FIC_0_AXI4_S_AWPROT({
        FIC_0_AXI4_S_AWPROT[2], FIC_0_AXI4_S_AWPROT[1], 
        FIC_0_AXI4_S_AWPROT[0]}), .FIC_0_AXI4_S_AWVALID(
        FIC_0_AXI4_S_AWVALID), .FIC_0_AXI4_S_WDATA({
        FIC_0_AXI4_S_WDATA[63], FIC_0_AXI4_S_WDATA[62], 
        FIC_0_AXI4_S_WDATA[61], FIC_0_AXI4_S_WDATA[60], 
        FIC_0_AXI4_S_WDATA[59], FIC_0_AXI4_S_WDATA[58], 
        FIC_0_AXI4_S_WDATA[57], FIC_0_AXI4_S_WDATA[56], 
        FIC_0_AXI4_S_WDATA[55], FIC_0_AXI4_S_WDATA[54], 
        FIC_0_AXI4_S_WDATA[53], FIC_0_AXI4_S_WDATA[52], 
        FIC_0_AXI4_S_WDATA[51], FIC_0_AXI4_S_WDATA[50], 
        FIC_0_AXI4_S_WDATA[49], FIC_0_AXI4_S_WDATA[48], 
        FIC_0_AXI4_S_WDATA[47], FIC_0_AXI4_S_WDATA[46], 
        FIC_0_AXI4_S_WDATA[45], FIC_0_AXI4_S_WDATA[44], 
        FIC_0_AXI4_S_WDATA[43], FIC_0_AXI4_S_WDATA[42], 
        FIC_0_AXI4_S_WDATA[41], FIC_0_AXI4_S_WDATA[40], 
        FIC_0_AXI4_S_WDATA[39], FIC_0_AXI4_S_WDATA[38], 
        FIC_0_AXI4_S_WDATA[37], FIC_0_AXI4_S_WDATA[36], 
        FIC_0_AXI4_S_WDATA[35], FIC_0_AXI4_S_WDATA[34], 
        FIC_0_AXI4_S_WDATA[33], FIC_0_AXI4_S_WDATA[32], 
        FIC_0_AXI4_S_WDATA[31], FIC_0_AXI4_S_WDATA[30], 
        FIC_0_AXI4_S_WDATA[29], FIC_0_AXI4_S_WDATA[28], 
        FIC_0_AXI4_S_WDATA[27], FIC_0_AXI4_S_WDATA[26], 
        FIC_0_AXI4_S_WDATA[25], FIC_0_AXI4_S_WDATA[24], 
        FIC_0_AXI4_S_WDATA[23], FIC_0_AXI4_S_WDATA[22], 
        FIC_0_AXI4_S_WDATA[21], FIC_0_AXI4_S_WDATA[20], 
        FIC_0_AXI4_S_WDATA[19], FIC_0_AXI4_S_WDATA[18], 
        FIC_0_AXI4_S_WDATA[17], FIC_0_AXI4_S_WDATA[16], 
        FIC_0_AXI4_S_WDATA[15], FIC_0_AXI4_S_WDATA[14], 
        FIC_0_AXI4_S_WDATA[13], FIC_0_AXI4_S_WDATA[12], 
        FIC_0_AXI4_S_WDATA[11], FIC_0_AXI4_S_WDATA[10], 
        FIC_0_AXI4_S_WDATA[9], FIC_0_AXI4_S_WDATA[8], 
        FIC_0_AXI4_S_WDATA[7], FIC_0_AXI4_S_WDATA[6], 
        FIC_0_AXI4_S_WDATA[5], FIC_0_AXI4_S_WDATA[4], 
        FIC_0_AXI4_S_WDATA[3], FIC_0_AXI4_S_WDATA[2], 
        FIC_0_AXI4_S_WDATA[1], FIC_0_AXI4_S_WDATA[0]}), 
        .FIC_0_AXI4_S_WSTRB({FIC_0_AXI4_S_WSTRB[7], 
        FIC_0_AXI4_S_WSTRB[6], FIC_0_AXI4_S_WSTRB[5], 
        FIC_0_AXI4_S_WSTRB[4], FIC_0_AXI4_S_WSTRB[3], 
        FIC_0_AXI4_S_WSTRB[2], FIC_0_AXI4_S_WSTRB[1], 
        FIC_0_AXI4_S_WSTRB[0]}), .FIC_0_AXI4_S_WLAST(
        FIC_0_AXI4_S_WLAST), .FIC_0_AXI4_S_WVALID(FIC_0_AXI4_S_WVALID), 
        .FIC_0_AXI4_S_BREADY(FIC_0_AXI4_S_BREADY), .FIC_0_AXI4_S_ARID({
        FIC_0_AXI4_S_ARID[3], FIC_0_AXI4_S_ARID[2], 
        FIC_0_AXI4_S_ARID[1], FIC_0_AXI4_S_ARID[0]}), 
        .FIC_0_AXI4_S_ARADDR({FIC_0_AXI4_S_ARADDR[37], 
        FIC_0_AXI4_S_ARADDR[36], FIC_0_AXI4_S_ARADDR[35], 
        FIC_0_AXI4_S_ARADDR[34], FIC_0_AXI4_S_ARADDR[33], 
        FIC_0_AXI4_S_ARADDR[32], FIC_0_AXI4_S_ARADDR[31], 
        FIC_0_AXI4_S_ARADDR[30], FIC_0_AXI4_S_ARADDR[29], 
        FIC_0_AXI4_S_ARADDR[28], FIC_0_AXI4_S_ARADDR[27], 
        FIC_0_AXI4_S_ARADDR[26], FIC_0_AXI4_S_ARADDR[25], 
        FIC_0_AXI4_S_ARADDR[24], FIC_0_AXI4_S_ARADDR[23], 
        FIC_0_AXI4_S_ARADDR[22], FIC_0_AXI4_S_ARADDR[21], 
        FIC_0_AXI4_S_ARADDR[20], FIC_0_AXI4_S_ARADDR[19], 
        FIC_0_AXI4_S_ARADDR[18], FIC_0_AXI4_S_ARADDR[17], 
        FIC_0_AXI4_S_ARADDR[16], FIC_0_AXI4_S_ARADDR[15], 
        FIC_0_AXI4_S_ARADDR[14], FIC_0_AXI4_S_ARADDR[13], 
        FIC_0_AXI4_S_ARADDR[12], FIC_0_AXI4_S_ARADDR[11], 
        FIC_0_AXI4_S_ARADDR[10], FIC_0_AXI4_S_ARADDR[9], 
        FIC_0_AXI4_S_ARADDR[8], FIC_0_AXI4_S_ARADDR[7], 
        FIC_0_AXI4_S_ARADDR[6], FIC_0_AXI4_S_ARADDR[5], 
        FIC_0_AXI4_S_ARADDR[4], FIC_0_AXI4_S_ARADDR[3], 
        FIC_0_AXI4_S_ARADDR[2], FIC_0_AXI4_S_ARADDR[1], 
        FIC_0_AXI4_S_ARADDR[0]}), .FIC_0_AXI4_S_ARLEN({
        FIC_0_AXI4_S_ARLEN[7], FIC_0_AXI4_S_ARLEN[6], 
        FIC_0_AXI4_S_ARLEN[5], FIC_0_AXI4_S_ARLEN[4], 
        FIC_0_AXI4_S_ARLEN[3], FIC_0_AXI4_S_ARLEN[2], 
        FIC_0_AXI4_S_ARLEN[1], FIC_0_AXI4_S_ARLEN[0]}), 
        .FIC_0_AXI4_S_ARSIZE({FIC_0_AXI4_S_ARSIZE[2], 
        FIC_0_AXI4_S_ARSIZE[1], FIC_0_AXI4_S_ARSIZE[0]}), 
        .FIC_0_AXI4_S_ARBURST({FIC_0_AXI4_S_ARBURST[1], 
        FIC_0_AXI4_S_ARBURST[0]}), .FIC_0_AXI4_S_ARQOS({
        FIC_0_AXI4_S_ARQOS[3], FIC_0_AXI4_S_ARQOS[2], 
        FIC_0_AXI4_S_ARQOS[1], FIC_0_AXI4_S_ARQOS[0]}), 
        .FIC_0_AXI4_S_ARLOCK(FIC_0_AXI4_S_ARLOCK), 
        .FIC_0_AXI4_S_ARCACHE({FIC_0_AXI4_S_ARCACHE[3], 
        FIC_0_AXI4_S_ARCACHE[2], FIC_0_AXI4_S_ARCACHE[1], 
        FIC_0_AXI4_S_ARCACHE[0]}), .FIC_0_AXI4_S_ARPROT({
        FIC_0_AXI4_S_ARPROT[2], FIC_0_AXI4_S_ARPROT[1], 
        FIC_0_AXI4_S_ARPROT[0]}), .FIC_0_AXI4_S_ARVALID(
        FIC_0_AXI4_S_ARVALID), .FIC_0_AXI4_S_RREADY(
        FIC_0_AXI4_S_RREADY), .FIC_1_ACLK(FIC_1_ACLK), 
        .FIC_1_AXI4_M_AWREADY(GND_net), .FIC_1_AXI4_M_WREADY(GND_net), 
        .FIC_1_AXI4_M_BID({GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net}), .FIC_1_AXI4_M_BRESP({GND_net, 
        GND_net}), .FIC_1_AXI4_M_BVALID(GND_net), 
        .FIC_1_AXI4_M_ARREADY(GND_net), .FIC_1_AXI4_M_RID({GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net})
        , .FIC_1_AXI4_M_RDATA({GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net}), .FIC_1_AXI4_M_RRESP({
        GND_net, GND_net}), .FIC_1_AXI4_M_RLAST(GND_net), 
        .FIC_1_AXI4_M_RVALID(GND_net), .FIC_1_AXI4_S_AWID({
        FIC_1_AXI4_S_AWID[3], FIC_1_AXI4_S_AWID[2], 
        FIC_1_AXI4_S_AWID[1], FIC_1_AXI4_S_AWID[0]}), 
        .FIC_1_AXI4_S_AWADDR({FIC_1_AXI4_S_AWADDR[37], 
        FIC_1_AXI4_S_AWADDR[36], FIC_1_AXI4_S_AWADDR[35], 
        FIC_1_AXI4_S_AWADDR[34], FIC_1_AXI4_S_AWADDR[33], 
        FIC_1_AXI4_S_AWADDR[32], FIC_1_AXI4_S_AWADDR[31], 
        FIC_1_AXI4_S_AWADDR[30], FIC_1_AXI4_S_AWADDR[29], 
        FIC_1_AXI4_S_AWADDR[28], FIC_1_AXI4_S_AWADDR[27], 
        FIC_1_AXI4_S_AWADDR[26], FIC_1_AXI4_S_AWADDR[25], 
        FIC_1_AXI4_S_AWADDR[24], FIC_1_AXI4_S_AWADDR[23], 
        FIC_1_AXI4_S_AWADDR[22], FIC_1_AXI4_S_AWADDR[21], 
        FIC_1_AXI4_S_AWADDR[20], FIC_1_AXI4_S_AWADDR[19], 
        FIC_1_AXI4_S_AWADDR[18], FIC_1_AXI4_S_AWADDR[17], 
        FIC_1_AXI4_S_AWADDR[16], FIC_1_AXI4_S_AWADDR[15], 
        FIC_1_AXI4_S_AWADDR[14], FIC_1_AXI4_S_AWADDR[13], 
        FIC_1_AXI4_S_AWADDR[12], FIC_1_AXI4_S_AWADDR[11], 
        FIC_1_AXI4_S_AWADDR[10], FIC_1_AXI4_S_AWADDR[9], 
        FIC_1_AXI4_S_AWADDR[8], FIC_1_AXI4_S_AWADDR[7], 
        FIC_1_AXI4_S_AWADDR[6], FIC_1_AXI4_S_AWADDR[5], 
        FIC_1_AXI4_S_AWADDR[4], FIC_1_AXI4_S_AWADDR[3], 
        FIC_1_AXI4_S_AWADDR[2], FIC_1_AXI4_S_AWADDR[1], 
        FIC_1_AXI4_S_AWADDR[0]}), .FIC_1_AXI4_S_AWLEN({
        FIC_1_AXI4_S_AWLEN[7], FIC_1_AXI4_S_AWLEN[6], 
        FIC_1_AXI4_S_AWLEN[5], FIC_1_AXI4_S_AWLEN[4], 
        FIC_1_AXI4_S_AWLEN[3], FIC_1_AXI4_S_AWLEN[2], 
        FIC_1_AXI4_S_AWLEN[1], FIC_1_AXI4_S_AWLEN[0]}), 
        .FIC_1_AXI4_S_AWSIZE({FIC_1_AXI4_S_AWSIZE[2], 
        FIC_1_AXI4_S_AWSIZE[1], FIC_1_AXI4_S_AWSIZE[0]}), 
        .FIC_1_AXI4_S_AWBURST({FIC_1_AXI4_S_AWBURST[1], 
        FIC_1_AXI4_S_AWBURST[0]}), .FIC_1_AXI4_S_AWLOCK(
        FIC_1_AXI4_S_AWLOCK), .FIC_1_AXI4_S_AWCACHE({
        FIC_1_AXI4_S_AWCACHE[3], FIC_1_AXI4_S_AWCACHE[2], 
        FIC_1_AXI4_S_AWCACHE[1], FIC_1_AXI4_S_AWCACHE[0]}), 
        .FIC_1_AXI4_S_AWQOS({FIC_1_AXI4_S_AWQOS[3], 
        FIC_1_AXI4_S_AWQOS[2], FIC_1_AXI4_S_AWQOS[1], 
        FIC_1_AXI4_S_AWQOS[0]}), .FIC_1_AXI4_S_AWPROT({
        FIC_1_AXI4_S_AWPROT[2], FIC_1_AXI4_S_AWPROT[1], 
        FIC_1_AXI4_S_AWPROT[0]}), .FIC_1_AXI4_S_AWVALID(
        FIC_1_AXI4_S_AWVALID), .FIC_1_AXI4_S_WDATA({
        FIC_1_AXI4_S_WDATA[63], FIC_1_AXI4_S_WDATA[62], 
        FIC_1_AXI4_S_WDATA[61], FIC_1_AXI4_S_WDATA[60], 
        FIC_1_AXI4_S_WDATA[59], FIC_1_AXI4_S_WDATA[58], 
        FIC_1_AXI4_S_WDATA[57], FIC_1_AXI4_S_WDATA[56], 
        FIC_1_AXI4_S_WDATA[55], FIC_1_AXI4_S_WDATA[54], 
        FIC_1_AXI4_S_WDATA[53], FIC_1_AXI4_S_WDATA[52], 
        FIC_1_AXI4_S_WDATA[51], FIC_1_AXI4_S_WDATA[50], 
        FIC_1_AXI4_S_WDATA[49], FIC_1_AXI4_S_WDATA[48], 
        FIC_1_AXI4_S_WDATA[47], FIC_1_AXI4_S_WDATA[46], 
        FIC_1_AXI4_S_WDATA[45], FIC_1_AXI4_S_WDATA[44], 
        FIC_1_AXI4_S_WDATA[43], FIC_1_AXI4_S_WDATA[42], 
        FIC_1_AXI4_S_WDATA[41], FIC_1_AXI4_S_WDATA[40], 
        FIC_1_AXI4_S_WDATA[39], FIC_1_AXI4_S_WDATA[38], 
        FIC_1_AXI4_S_WDATA[37], FIC_1_AXI4_S_WDATA[36], 
        FIC_1_AXI4_S_WDATA[35], FIC_1_AXI4_S_WDATA[34], 
        FIC_1_AXI4_S_WDATA[33], FIC_1_AXI4_S_WDATA[32], 
        FIC_1_AXI4_S_WDATA[31], FIC_1_AXI4_S_WDATA[30], 
        FIC_1_AXI4_S_WDATA[29], FIC_1_AXI4_S_WDATA[28], 
        FIC_1_AXI4_S_WDATA[27], FIC_1_AXI4_S_WDATA[26], 
        FIC_1_AXI4_S_WDATA[25], FIC_1_AXI4_S_WDATA[24], 
        FIC_1_AXI4_S_WDATA[23], FIC_1_AXI4_S_WDATA[22], 
        FIC_1_AXI4_S_WDATA[21], FIC_1_AXI4_S_WDATA[20], 
        FIC_1_AXI4_S_WDATA[19], FIC_1_AXI4_S_WDATA[18], 
        FIC_1_AXI4_S_WDATA[17], FIC_1_AXI4_S_WDATA[16], 
        FIC_1_AXI4_S_WDATA[15], FIC_1_AXI4_S_WDATA[14], 
        FIC_1_AXI4_S_WDATA[13], FIC_1_AXI4_S_WDATA[12], 
        FIC_1_AXI4_S_WDATA[11], FIC_1_AXI4_S_WDATA[10], 
        FIC_1_AXI4_S_WDATA[9], FIC_1_AXI4_S_WDATA[8], 
        FIC_1_AXI4_S_WDATA[7], FIC_1_AXI4_S_WDATA[6], 
        FIC_1_AXI4_S_WDATA[5], FIC_1_AXI4_S_WDATA[4], 
        FIC_1_AXI4_S_WDATA[3], FIC_1_AXI4_S_WDATA[2], 
        FIC_1_AXI4_S_WDATA[1], FIC_1_AXI4_S_WDATA[0]}), 
        .FIC_1_AXI4_S_WSTRB({FIC_1_AXI4_S_WSTRB[7], 
        FIC_1_AXI4_S_WSTRB[6], FIC_1_AXI4_S_WSTRB[5], 
        FIC_1_AXI4_S_WSTRB[4], FIC_1_AXI4_S_WSTRB[3], 
        FIC_1_AXI4_S_WSTRB[2], FIC_1_AXI4_S_WSTRB[1], 
        FIC_1_AXI4_S_WSTRB[0]}), .FIC_1_AXI4_S_WLAST(
        FIC_1_AXI4_S_WLAST), .FIC_1_AXI4_S_WVALID(FIC_1_AXI4_S_WVALID), 
        .FIC_1_AXI4_S_BREADY(FIC_1_AXI4_S_BREADY), .FIC_1_AXI4_S_ARID({
        FIC_1_AXI4_S_ARID[3], FIC_1_AXI4_S_ARID[2], 
        FIC_1_AXI4_S_ARID[1], FIC_1_AXI4_S_ARID[0]}), 
        .FIC_1_AXI4_S_ARADDR({FIC_1_AXI4_S_ARADDR[37], 
        FIC_1_AXI4_S_ARADDR[36], FIC_1_AXI4_S_ARADDR[35], 
        FIC_1_AXI4_S_ARADDR[34], FIC_1_AXI4_S_ARADDR[33], 
        FIC_1_AXI4_S_ARADDR[32], FIC_1_AXI4_S_ARADDR[31], 
        FIC_1_AXI4_S_ARADDR[30], FIC_1_AXI4_S_ARADDR[29], 
        FIC_1_AXI4_S_ARADDR[28], FIC_1_AXI4_S_ARADDR[27], 
        FIC_1_AXI4_S_ARADDR[26], FIC_1_AXI4_S_ARADDR[25], 
        FIC_1_AXI4_S_ARADDR[24], FIC_1_AXI4_S_ARADDR[23], 
        FIC_1_AXI4_S_ARADDR[22], FIC_1_AXI4_S_ARADDR[21], 
        FIC_1_AXI4_S_ARADDR[20], FIC_1_AXI4_S_ARADDR[19], 
        FIC_1_AXI4_S_ARADDR[18], FIC_1_AXI4_S_ARADDR[17], 
        FIC_1_AXI4_S_ARADDR[16], FIC_1_AXI4_S_ARADDR[15], 
        FIC_1_AXI4_S_ARADDR[14], FIC_1_AXI4_S_ARADDR[13], 
        FIC_1_AXI4_S_ARADDR[12], FIC_1_AXI4_S_ARADDR[11], 
        FIC_1_AXI4_S_ARADDR[10], FIC_1_AXI4_S_ARADDR[9], 
        FIC_1_AXI4_S_ARADDR[8], FIC_1_AXI4_S_ARADDR[7], 
        FIC_1_AXI4_S_ARADDR[6], FIC_1_AXI4_S_ARADDR[5], 
        FIC_1_AXI4_S_ARADDR[4], FIC_1_AXI4_S_ARADDR[3], 
        FIC_1_AXI4_S_ARADDR[2], FIC_1_AXI4_S_ARADDR[1], 
        FIC_1_AXI4_S_ARADDR[0]}), .FIC_1_AXI4_S_ARLEN({
        FIC_1_AXI4_S_ARLEN[7], FIC_1_AXI4_S_ARLEN[6], 
        FIC_1_AXI4_S_ARLEN[5], FIC_1_AXI4_S_ARLEN[4], 
        FIC_1_AXI4_S_ARLEN[3], FIC_1_AXI4_S_ARLEN[2], 
        FIC_1_AXI4_S_ARLEN[1], FIC_1_AXI4_S_ARLEN[0]}), 
        .FIC_1_AXI4_S_ARSIZE({FIC_1_AXI4_S_ARSIZE[2], 
        FIC_1_AXI4_S_ARSIZE[1], FIC_1_AXI4_S_ARSIZE[0]}), 
        .FIC_1_AXI4_S_ARBURST({FIC_1_AXI4_S_ARBURST[1], 
        FIC_1_AXI4_S_ARBURST[0]}), .FIC_1_AXI4_S_ARQOS({
        FIC_1_AXI4_S_ARQOS[3], FIC_1_AXI4_S_ARQOS[2], 
        FIC_1_AXI4_S_ARQOS[1], FIC_1_AXI4_S_ARQOS[0]}), 
        .FIC_1_AXI4_S_ARLOCK(FIC_1_AXI4_S_ARLOCK), 
        .FIC_1_AXI4_S_ARCACHE({FIC_1_AXI4_S_ARCACHE[3], 
        FIC_1_AXI4_S_ARCACHE[2], FIC_1_AXI4_S_ARCACHE[1], 
        FIC_1_AXI4_S_ARCACHE[0]}), .FIC_1_AXI4_S_ARPROT({
        FIC_1_AXI4_S_ARPROT[2], FIC_1_AXI4_S_ARPROT[1], 
        FIC_1_AXI4_S_ARPROT[0]}), .FIC_1_AXI4_S_ARVALID(
        FIC_1_AXI4_S_ARVALID), .FIC_1_AXI4_S_RREADY(
        FIC_1_AXI4_S_RREADY), .FIC_2_ACLK(FIC_2_ACLK), .SPARE_3_F2M(
        FIC_3_APB_M_PADDR[30]), .FIC_2_AXI4_S_AWID({
        FIC_2_AXI4_S_AWID[3], FIC_2_AXI4_S_AWID[2], 
        FIC_2_AXI4_S_AWID[1], FIC_2_AXI4_S_AWID[0]}), 
        .FIC_2_AXI4_S_AWADDR({FIC_2_AXI4_S_AWADDR[37], 
        FIC_2_AXI4_S_AWADDR[36], FIC_2_AXI4_S_AWADDR[35], 
        FIC_2_AXI4_S_AWADDR[34], FIC_2_AXI4_S_AWADDR[33], 
        FIC_2_AXI4_S_AWADDR[32], FIC_2_AXI4_S_AWADDR[31], 
        FIC_2_AXI4_S_AWADDR[30], FIC_2_AXI4_S_AWADDR[29], 
        FIC_2_AXI4_S_AWADDR[28], FIC_2_AXI4_S_AWADDR[27], 
        FIC_2_AXI4_S_AWADDR[26], FIC_2_AXI4_S_AWADDR[25], 
        FIC_2_AXI4_S_AWADDR[24], FIC_2_AXI4_S_AWADDR[23], 
        FIC_2_AXI4_S_AWADDR[22], FIC_2_AXI4_S_AWADDR[21], 
        FIC_2_AXI4_S_AWADDR[20], FIC_2_AXI4_S_AWADDR[19], 
        FIC_2_AXI4_S_AWADDR[18], FIC_2_AXI4_S_AWADDR[17], 
        FIC_2_AXI4_S_AWADDR[16], FIC_2_AXI4_S_AWADDR[15], 
        FIC_2_AXI4_S_AWADDR[14], FIC_2_AXI4_S_AWADDR[13], 
        FIC_2_AXI4_S_AWADDR[12], FIC_2_AXI4_S_AWADDR[11], 
        FIC_2_AXI4_S_AWADDR[10], FIC_2_AXI4_S_AWADDR[9], 
        FIC_2_AXI4_S_AWADDR[8], FIC_2_AXI4_S_AWADDR[7], 
        FIC_2_AXI4_S_AWADDR[6], FIC_2_AXI4_S_AWADDR[5], 
        FIC_2_AXI4_S_AWADDR[4], FIC_2_AXI4_S_AWADDR[3], 
        FIC_2_AXI4_S_AWADDR[2], FIC_2_AXI4_S_AWADDR[1], 
        FIC_2_AXI4_S_AWADDR[0]}), .FIC_2_AXI4_S_AWLEN({
        FIC_2_AXI4_S_AWLEN[7], FIC_2_AXI4_S_AWLEN[6], 
        FIC_2_AXI4_S_AWLEN[5], FIC_2_AXI4_S_AWLEN[4], 
        FIC_2_AXI4_S_AWLEN[3], FIC_2_AXI4_S_AWLEN[2], 
        FIC_2_AXI4_S_AWLEN[1], FIC_2_AXI4_S_AWLEN[0]}), 
        .FIC_2_AXI4_S_AWSIZE({FIC_2_AXI4_S_AWSIZE[2], 
        FIC_2_AXI4_S_AWSIZE[1], FIC_2_AXI4_S_AWSIZE[0]}), 
        .FIC_2_AXI4_S_AWBURST({FIC_2_AXI4_S_AWBURST[1], 
        FIC_2_AXI4_S_AWBURST[0]}), .FIC_2_AXI4_S_AWLOCK(
        FIC_2_AXI4_S_AWLOCK), .FIC_2_AXI4_S_AWCACHE({
        FIC_2_AXI4_S_AWCACHE[3], FIC_2_AXI4_S_AWCACHE[2], 
        FIC_2_AXI4_S_AWCACHE[1], FIC_2_AXI4_S_AWCACHE[0]}), 
        .FIC_2_AXI4_S_AWQOS({FIC_2_AXI4_S_AWQOS[3], 
        FIC_2_AXI4_S_AWQOS[2], FIC_2_AXI4_S_AWQOS[1], 
        FIC_2_AXI4_S_AWQOS[0]}), .FIC_2_AXI4_S_AWPROT({
        FIC_2_AXI4_S_AWPROT[2], FIC_2_AXI4_S_AWPROT[1], 
        FIC_2_AXI4_S_AWPROT[0]}), .FIC_2_AXI4_S_AWVALID(
        FIC_2_AXI4_S_AWVALID), .FIC_2_AXI4_S_WDATA({
        FIC_2_AXI4_S_WDATA[63], FIC_2_AXI4_S_WDATA[62], 
        FIC_2_AXI4_S_WDATA[61], FIC_2_AXI4_S_WDATA[60], 
        FIC_2_AXI4_S_WDATA[59], FIC_2_AXI4_S_WDATA[58], 
        FIC_2_AXI4_S_WDATA[57], FIC_2_AXI4_S_WDATA[56], 
        FIC_2_AXI4_S_WDATA[55], FIC_2_AXI4_S_WDATA[54], 
        FIC_2_AXI4_S_WDATA[53], FIC_2_AXI4_S_WDATA[52], 
        FIC_2_AXI4_S_WDATA[51], FIC_2_AXI4_S_WDATA[50], 
        FIC_2_AXI4_S_WDATA[49], FIC_2_AXI4_S_WDATA[48], 
        FIC_2_AXI4_S_WDATA[47], FIC_2_AXI4_S_WDATA[46], 
        FIC_2_AXI4_S_WDATA[45], FIC_2_AXI4_S_WDATA[44], 
        FIC_2_AXI4_S_WDATA[43], FIC_2_AXI4_S_WDATA[42], 
        FIC_2_AXI4_S_WDATA[41], FIC_2_AXI4_S_WDATA[40], 
        FIC_2_AXI4_S_WDATA[39], FIC_2_AXI4_S_WDATA[38], 
        FIC_2_AXI4_S_WDATA[37], FIC_2_AXI4_S_WDATA[36], 
        FIC_2_AXI4_S_WDATA[35], FIC_2_AXI4_S_WDATA[34], 
        FIC_2_AXI4_S_WDATA[33], FIC_2_AXI4_S_WDATA[32], 
        FIC_2_AXI4_S_WDATA[31], FIC_2_AXI4_S_WDATA[30], 
        FIC_2_AXI4_S_WDATA[29], FIC_2_AXI4_S_WDATA[28], 
        FIC_2_AXI4_S_WDATA[27], FIC_2_AXI4_S_WDATA[26], 
        FIC_2_AXI4_S_WDATA[25], FIC_2_AXI4_S_WDATA[24], 
        FIC_2_AXI4_S_WDATA[23], FIC_2_AXI4_S_WDATA[22], 
        FIC_2_AXI4_S_WDATA[21], FIC_2_AXI4_S_WDATA[20], 
        FIC_2_AXI4_S_WDATA[19], FIC_2_AXI4_S_WDATA[18], 
        FIC_2_AXI4_S_WDATA[17], FIC_2_AXI4_S_WDATA[16], 
        FIC_2_AXI4_S_WDATA[15], FIC_2_AXI4_S_WDATA[14], 
        FIC_2_AXI4_S_WDATA[13], FIC_2_AXI4_S_WDATA[12], 
        FIC_2_AXI4_S_WDATA[11], FIC_2_AXI4_S_WDATA[10], 
        FIC_2_AXI4_S_WDATA[9], FIC_2_AXI4_S_WDATA[8], 
        FIC_2_AXI4_S_WDATA[7], FIC_2_AXI4_S_WDATA[6], 
        FIC_2_AXI4_S_WDATA[5], FIC_2_AXI4_S_WDATA[4], 
        FIC_2_AXI4_S_WDATA[3], FIC_2_AXI4_S_WDATA[2], 
        FIC_2_AXI4_S_WDATA[1], FIC_2_AXI4_S_WDATA[0]}), 
        .FIC_2_AXI4_S_WSTRB({FIC_2_AXI4_S_WSTRB[7], 
        FIC_2_AXI4_S_WSTRB[6], FIC_2_AXI4_S_WSTRB[5], 
        FIC_2_AXI4_S_WSTRB[4], FIC_2_AXI4_S_WSTRB[3], 
        FIC_2_AXI4_S_WSTRB[2], FIC_2_AXI4_S_WSTRB[1], 
        FIC_2_AXI4_S_WSTRB[0]}), .FIC_2_AXI4_S_WLAST(
        FIC_2_AXI4_S_WLAST), .FIC_2_AXI4_S_WVALID(FIC_2_AXI4_S_WVALID), 
        .FIC_2_AXI4_S_BREADY(FIC_2_AXI4_S_BREADY), .FIC_2_AXI4_S_ARID({
        FIC_2_AXI4_S_ARID[3], FIC_2_AXI4_S_ARID[2], 
        FIC_2_AXI4_S_ARID[1], FIC_2_AXI4_S_ARID[0]}), 
        .FIC_2_AXI4_S_ARADDR({FIC_2_AXI4_S_ARADDR[37], 
        FIC_2_AXI4_S_ARADDR[36], FIC_2_AXI4_S_ARADDR[35], 
        FIC_2_AXI4_S_ARADDR[34], FIC_2_AXI4_S_ARADDR[33], 
        FIC_2_AXI4_S_ARADDR[32], FIC_2_AXI4_S_ARADDR[31], 
        FIC_2_AXI4_S_ARADDR[30], FIC_2_AXI4_S_ARADDR[29], 
        FIC_2_AXI4_S_ARADDR[28], FIC_2_AXI4_S_ARADDR[27], 
        FIC_2_AXI4_S_ARADDR[26], FIC_2_AXI4_S_ARADDR[25], 
        FIC_2_AXI4_S_ARADDR[24], FIC_2_AXI4_S_ARADDR[23], 
        FIC_2_AXI4_S_ARADDR[22], FIC_2_AXI4_S_ARADDR[21], 
        FIC_2_AXI4_S_ARADDR[20], FIC_2_AXI4_S_ARADDR[19], 
        FIC_2_AXI4_S_ARADDR[18], FIC_2_AXI4_S_ARADDR[17], 
        FIC_2_AXI4_S_ARADDR[16], FIC_2_AXI4_S_ARADDR[15], 
        FIC_2_AXI4_S_ARADDR[14], FIC_2_AXI4_S_ARADDR[13], 
        FIC_2_AXI4_S_ARADDR[12], FIC_2_AXI4_S_ARADDR[11], 
        FIC_2_AXI4_S_ARADDR[10], FIC_2_AXI4_S_ARADDR[9], 
        FIC_2_AXI4_S_ARADDR[8], FIC_2_AXI4_S_ARADDR[7], 
        FIC_2_AXI4_S_ARADDR[6], FIC_2_AXI4_S_ARADDR[5], 
        FIC_2_AXI4_S_ARADDR[4], FIC_2_AXI4_S_ARADDR[3], 
        FIC_2_AXI4_S_ARADDR[2], FIC_2_AXI4_S_ARADDR[1], 
        FIC_2_AXI4_S_ARADDR[0]}), .FIC_2_AXI4_S_ARLEN({
        FIC_2_AXI4_S_ARLEN[7], FIC_2_AXI4_S_ARLEN[6], 
        FIC_2_AXI4_S_ARLEN[5], FIC_2_AXI4_S_ARLEN[4], 
        FIC_2_AXI4_S_ARLEN[3], FIC_2_AXI4_S_ARLEN[2], 
        FIC_2_AXI4_S_ARLEN[1], FIC_2_AXI4_S_ARLEN[0]}), 
        .FIC_2_AXI4_S_ARSIZE({FIC_2_AXI4_S_ARSIZE[2], 
        FIC_2_AXI4_S_ARSIZE[1], FIC_2_AXI4_S_ARSIZE[0]}), 
        .FIC_2_AXI4_S_ARBURST({FIC_2_AXI4_S_ARBURST[1], 
        FIC_2_AXI4_S_ARBURST[0]}), .FIC_2_AXI4_S_ARLOCK(
        FIC_2_AXI4_S_ARLOCK), .FIC_2_AXI4_S_ARCACHE({
        FIC_2_AXI4_S_ARCACHE[3], FIC_2_AXI4_S_ARCACHE[2], 
        FIC_2_AXI4_S_ARCACHE[1], FIC_2_AXI4_S_ARCACHE[0]}), 
        .FIC_2_AXI4_S_ARQOS({FIC_2_AXI4_S_ARQOS[3], 
        FIC_2_AXI4_S_ARQOS[2], FIC_2_AXI4_S_ARQOS[1], 
        FIC_2_AXI4_S_ARQOS[0]}), .FIC_2_AXI4_S_ARPROT({
        FIC_2_AXI4_S_ARPROT[2], FIC_2_AXI4_S_ARPROT[1], 
        FIC_2_AXI4_S_ARPROT[0]}), .FIC_2_AXI4_S_ARVALID(
        FIC_2_AXI4_S_ARVALID), .FIC_2_AXI4_S_RREADY(
        FIC_2_AXI4_S_RREADY), .FIC_3_PCLK(FIC_3_PCLK), .SPARE_4_F2M(
        FIC_3_APB_M_PADDR[30]), .FIC_3_APB_M_PRDATA({
        FIC_3_APB_M_PRDATA[31], FIC_3_APB_M_PRDATA[30], 
        FIC_3_APB_M_PRDATA[29], FIC_3_APB_M_PRDATA[28], 
        FIC_3_APB_M_PRDATA[27], FIC_3_APB_M_PRDATA[26], 
        FIC_3_APB_M_PRDATA[25], FIC_3_APB_M_PRDATA[24], 
        FIC_3_APB_M_PRDATA[23], FIC_3_APB_M_PRDATA[22], 
        FIC_3_APB_M_PRDATA[21], FIC_3_APB_M_PRDATA[20], 
        FIC_3_APB_M_PRDATA[19], FIC_3_APB_M_PRDATA[18], 
        FIC_3_APB_M_PRDATA[17], FIC_3_APB_M_PRDATA[16], 
        FIC_3_APB_M_PRDATA[15], FIC_3_APB_M_PRDATA[14], 
        FIC_3_APB_M_PRDATA[13], FIC_3_APB_M_PRDATA[12], 
        FIC_3_APB_M_PRDATA[11], FIC_3_APB_M_PRDATA[10], 
        FIC_3_APB_M_PRDATA[9], FIC_3_APB_M_PRDATA[8], 
        FIC_3_APB_M_PRDATA[7], FIC_3_APB_M_PRDATA[6], 
        FIC_3_APB_M_PRDATA[5], FIC_3_APB_M_PRDATA[4], 
        FIC_3_APB_M_PRDATA[3], FIC_3_APB_M_PRDATA[2], 
        FIC_3_APB_M_PRDATA[1], FIC_3_APB_M_PRDATA[0]}), 
        .FIC_3_APB_M_PREADY(FIC_3_APB_M_PREADY), .FIC_3_APB_M_PSLVERR(
        FIC_3_APB_M_PSLVERR), .MMUART_0_DCD_F2M(GND_net), 
        .MMUART_0_RI_F2M(GND_net), .MMUART_0_DSR_F2M(GND_net), 
        .MMUART_0_CTS_F2M(GND_net), .MMUART_0_RXD_F2M(MMUART_0_RXD_F2M)
        , .MMUART_0_CLK_F2M(GND_net), .MMUART_1_DCD_F2M(GND_net), 
        .MMUART_1_RI_F2M(GND_net), .MMUART_1_DSR_F2M(GND_net), 
        .MMUART_1_CTS_F2M(GND_net), .MMUART_1_RXD_F2M(MMUART_1_RXD_F2M)
        , .MMUART_1_CLK_F2M(GND_net), .MMUART_2_RXD_F2M(
        MMUART_2_RXD_F2M), .MMUART_3_RXD_F2M(MMUART_3_RXD_F2M), 
        .MMUART_4_RXD_F2M(MMUART_4_RXD_F2M), .CAN_0_RXBUS_F2M(
        CAN_0_RXBUS_F2M), .CAN_1_RXBUS_F2M(GND_net), .CAN_CLK_F2M(
        FIC_3_APB_M_PADDR[30]), .QSPI_DATA_F2M({QSPI_DATA3_F2M, 
        QSPI_DATA2_F2M, GND_net, GND_net}), .SPI_0_SS_F2M(SPI_0_SS_F2M)
        , .SPI_0_DI_F2M(SPI_0_DI_F2M), .SPI_0_CLK_F2M(SPI_0_CLK_F2M), 
        .SPI_1_SS_F2M(GND_net), .SPI_1_DI_F2M(GND_net), .SPI_1_CLK_F2M(
        GND_net), .I2C_0_SCL_F2M(I2C_0_SCL_F2M), .I2C_1_SCL_F2M(
        GND_net), .I2C_0_SDA_F2M(I2C_0_SDA_F2M), .I2C_1_SDA_F2M(
        GND_net), .I2C_0_BCLK_F2M(GND_net), .I2C_0_SMBALERT_NI_F2M(
        GND_net), .I2C_0_SMBSUS_NI_F2M(GND_net), .I2C_1_BCLK_F2M(
        GND_net), .I2C_1_SMBALERT_NI_F2M(GND_net), 
        .I2C_1_SMBSUS_NI_F2M(GND_net), .GPIO_2_F2M({GPIO_2_F2M_31, 
        GPIO_2_F2M_30, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net}), .MAC_0_MDI_F2M(GND_net), 
        .MAC_1_MDI_F2M(GND_net), .JTAG_TMS_F2M(GND_net), .JTAG_TCK_F2M(
        GND_net), .JTAG_TDI_F2M(GND_net), .JTAG_TRSTB_F2M(GND_net), 
        .MSS_INT_F2M({MSS_INT_F2M[63], MSS_INT_F2M[62], 
        MSS_INT_F2M[61], MSS_INT_F2M[60], MSS_INT_F2M[59], 
        MSS_INT_F2M[58], MSS_INT_F2M[57], MSS_INT_F2M[56], 
        MSS_INT_F2M[55], MSS_INT_F2M[54], MSS_INT_F2M[53], 
        MSS_INT_F2M[52], MSS_INT_F2M[51], MSS_INT_F2M[50], 
        MSS_INT_F2M[49], MSS_INT_F2M[48], MSS_INT_F2M[47], 
        MSS_INT_F2M[46], MSS_INT_F2M[45], MSS_INT_F2M[44], 
        MSS_INT_F2M[43], MSS_INT_F2M[42], MSS_INT_F2M[41], 
        MSS_INT_F2M[40], MSS_INT_F2M[39], MSS_INT_F2M[38], 
        MSS_INT_F2M[37], MSS_INT_F2M[36], MSS_INT_F2M[35], 
        MSS_INT_F2M[34], MSS_INT_F2M[33], MSS_INT_F2M[32], 
        MSS_INT_F2M[31], MSS_INT_F2M[30], MSS_INT_F2M[29], 
        MSS_INT_F2M[28], MSS_INT_F2M[27], MSS_INT_F2M[26], 
        MSS_INT_F2M[25], MSS_INT_F2M[24], MSS_INT_F2M[23], 
        MSS_INT_F2M[22], MSS_INT_F2M[21], MSS_INT_F2M[20], 
        MSS_INT_F2M[19], MSS_INT_F2M[18], MSS_INT_F2M[17], 
        MSS_INT_F2M[16], MSS_INT_F2M[15], MSS_INT_F2M[14], 
        MSS_INT_F2M[13], MSS_INT_F2M[12], MSS_INT_F2M[11], 
        MSS_INT_F2M[10], MSS_INT_F2M[9], MSS_INT_F2M[8], 
        MSS_INT_F2M[7], MSS_INT_F2M[6], MSS_INT_F2M[5], MSS_INT_F2M[4], 
        MSS_INT_F2M[3], MSS_INT_F2M[2], MSS_INT_F2M[1], MSS_INT_F2M[0]})
        , .SPARE_1_F2M({GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net}), .SPARE_2_F2M({
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net}), .BOOT_FAIL_CLEAR_F2M(GND_net), 
        .MSS_RESET_N_F2M(MSS_RESET_N_F2M), .GPIO_RESET_N_F2M(GND_net), 
        .USOC_TRACE_CLOCK_F2M(GND_net), .USOC_TRACE_VALID_F2M(GND_net), 
        .USOC_TRACE_DATA_F2M({GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net}), .SPARE_5_F2M(FIC_3_APB_M_PADDR[30]), 
        .MAC_0_GMII_MII_RXD_F2M({GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net}), 
        .MAC_0_GMII_MII_RX_DV_F2M(GND_net), .MAC_0_GMII_MII_RX_ER_F2M(
        GND_net), .MAC_0_GMII_MII_RX_CRS_F2M(GND_net), 
        .MAC_0_GMII_MII_RX_COL_F2M(GND_net), 
        .MAC_0_GMII_MII_RX_CLK_F2M(GND_net), 
        .MAC_0_GMII_MII_TX_CLK_F2M(GND_net), .MAC_0_TSU_CLK_F2M(
        GND_net), .MAC_1_GMII_MII_RXD_F2M({GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net}), 
        .MAC_1_GMII_MII_RX_DV_F2M(GND_net), .MAC_1_GMII_MII_RX_ER_F2M(
        GND_net), .MAC_1_GMII_MII_RX_CRS_F2M(GND_net), 
        .MAC_1_GMII_MII_RX_COL_F2M(GND_net), 
        .MAC_1_GMII_MII_RX_CLK_F2M(GND_net), 
        .MAC_1_GMII_MII_TX_CLK_F2M(GND_net), .MAC_1_TSU_CLK_F2M(
        GND_net), .MAC_0_FILTER_MATCH1_F2M(GND_net), 
        .MAC_0_FILTER_MATCH2_F2M(GND_net), .MAC_0_FILTER_MATCH3_F2M(
        GND_net), .MAC_0_FILTER_MATCH4_F2M(GND_net), 
        .MAC_1_FILTER_MATCH1_F2M(GND_net), .MAC_1_FILTER_MATCH2_F2M(
        GND_net), .MAC_1_FILTER_MATCH3_F2M(GND_net), 
        .MAC_1_FILTER_MATCH4_F2M(GND_net), .MAC_0_TSU_GEM_MS_F2M(
        GND_net), .MAC_0_TSU_GEM_INC_CTRL_F2M({GND_net, GND_net}), 
        .MAC_1_TSU_GEM_MS_F2M(GND_net), .MAC_1_TSU_GEM_INC_CTRL_F2M({
        GND_net, GND_net}), .CRYPTO_HCLK(FIC_3_APB_M_PADDR[30]), 
        .CRYPTO_HRESETN(FIC_3_APB_M_PADDR[30]), .CRYPTO_AHB_M_HREADY(
        GND_net), .CRYPTO_AHB_M_HRESP(GND_net), .CRYPTO_AHB_M_HRDATA({
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net}), .CRYPTO_AHB_S_HSEL(
        GND_net), .CRYPTO_AHB_S_HADDR({GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net})
        , .CRYPTO_AHB_S_HWDATA({GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net})
        , .CRYPTO_AHB_S_HSIZE({GND_net, GND_net}), 
        .CRYPTO_AHB_S_HTRANS({GND_net, GND_net}), .CRYPTO_AHB_S_HWRITE(
        GND_net), .CRYPTO_AHB_S_HREADY(GND_net), .CRYPTO_STALL_F2M(
        FIC_3_APB_M_PADDR[30]), .CRYPTO_PURGE_F2M(
        FIC_3_APB_M_PADDR[30]), .CRYPTO_GO_F2M(FIC_3_APB_M_PADDR[30]), 
        .CRYPTO_REQUEST_F2M(FIC_3_APB_M_PADDR[30]), 
        .CRYPTO_RELEASE_F2M(FIC_3_APB_M_PADDR[30]), 
        .CRYPTO_XENABLE_F2M(FIC_3_APB_M_PADDR[30]), .CRYPTO_XWDATA_F2M({
        FIC_3_APB_M_PADDR[30], FIC_3_APB_M_PADDR[30], 
        FIC_3_APB_M_PADDR[30], FIC_3_APB_M_PADDR[30], 
        FIC_3_APB_M_PADDR[30], FIC_3_APB_M_PADDR[30], 
        FIC_3_APB_M_PADDR[30], FIC_3_APB_M_PADDR[30], 
        FIC_3_APB_M_PADDR[30], FIC_3_APB_M_PADDR[30], 
        FIC_3_APB_M_PADDR[30], FIC_3_APB_M_PADDR[30], 
        FIC_3_APB_M_PADDR[30], FIC_3_APB_M_PADDR[30], 
        FIC_3_APB_M_PADDR[30], FIC_3_APB_M_PADDR[30], 
        FIC_3_APB_M_PADDR[30], FIC_3_APB_M_PADDR[30], 
        FIC_3_APB_M_PADDR[30], FIC_3_APB_M_PADDR[30], 
        FIC_3_APB_M_PADDR[30], FIC_3_APB_M_PADDR[30], 
        FIC_3_APB_M_PADDR[30], FIC_3_APB_M_PADDR[30], 
        FIC_3_APB_M_PADDR[30], FIC_3_APB_M_PADDR[30], 
        FIC_3_APB_M_PADDR[30], FIC_3_APB_M_PADDR[30], 
        FIC_3_APB_M_PADDR[30], FIC_3_APB_M_PADDR[30], 
        FIC_3_APB_M_PADDR[30], FIC_3_APB_M_PADDR[30]}), 
        .CRYPTO_XOUTACK_F2M(FIC_3_APB_M_PADDR[30]), 
        .CRYPTO_MESH_CLEAR_F2M(GND_net), .EMMC_SD_CLK_F2M(
        FIC_3_APB_M_PADDR[30]), .MSSIO37_IN(GND_net), .MSSIO37_OUT(), 
        .MSSIO37_OE(), .MSSIO36_IN(GND_net), .MSSIO36_OUT(
        D_MSSIO36_OUT_IOINST_net), .MSSIO36_OE(), .MSSIO35_IN(
        Y_MSSIO35_IN_IOINST_net), .MSSIO35_OUT(), .MSSIO35_OE(), 
        .MSSIO34_IN(GND_net), .MSSIO34_OUT(D_MSSIO34_OUT_IOINST_net), 
        .MSSIO34_OE(), .MSSIO33_IN(Y_MSSIO33_OUT_IOINST_net), 
        .MSSIO33_OUT(D_MSSIO33_OUT_IOINST_net), .MSSIO33_OE(
        E_MSSIO33_OUT_IOINST_net), .MSSIO32_IN(
        Y_MSSIO32_OUT_IOINST_net), .MSSIO32_OUT(
        D_MSSIO32_OUT_IOINST_net), .MSSIO32_OE(
        E_MSSIO32_OUT_IOINST_net), .MSSIO31_IN(GND_net), .MSSIO31_OUT(
        D_MSSIO31_OUT_IOINST_net), .MSSIO31_OE(), .MSSIO30_IN(GND_net), 
        .MSSIO30_OUT(D_MSSIO30_OUT_IOINST_net), .MSSIO30_OE(), 
        .MSSIO29_IN(Y_MSSIO29_OUT_IOINST_net), .MSSIO29_OUT(
        D_MSSIO29_OUT_IOINST_net), .MSSIO29_OE(
        E_MSSIO29_OUT_IOINST_net), .MSSIO28_IN(GND_net), .MSSIO28_OUT(
        D_MSSIO28_OUT_IOINST_net), .MSSIO28_OE(), .MSSIO27_IN(
        Y_MSSIO27_OUT_IOINST_net), .MSSIO27_OUT(
        D_MSSIO27_OUT_IOINST_net), .MSSIO27_OE(
        E_MSSIO27_OUT_IOINST_net), .MSSIO26_IN(
        Y_MSSIO26_OUT_IOINST_net), .MSSIO26_OUT(
        D_MSSIO26_OUT_IOINST_net), .MSSIO26_OE(
        E_MSSIO26_OUT_IOINST_net), .MSSIO25_IN(
        Y_MSSIO25_OUT_IOINST_net), .MSSIO25_OUT(
        D_MSSIO25_OUT_IOINST_net), .MSSIO25_OE(
        E_MSSIO25_OUT_IOINST_net), .MSSIO24_IN(
        Y_MSSIO24_OUT_IOINST_net), .MSSIO24_OUT(
        D_MSSIO24_OUT_IOINST_net), .MSSIO24_OE(
        E_MSSIO24_OUT_IOINST_net), .MSSIO23_IN(
        Y_MSSIO23_OUT_IOINST_net), .MSSIO23_OUT(
        D_MSSIO23_OUT_IOINST_net), .MSSIO23_OE(
        E_MSSIO23_OUT_IOINST_net), .MSSIO22_IN(
        Y_MSSIO22_OUT_IOINST_net), .MSSIO22_OUT(
        D_MSSIO22_OUT_IOINST_net), .MSSIO22_OE(
        E_MSSIO22_OUT_IOINST_net), .MSSIO21_IN(
        Y_MSSIO21_OUT_IOINST_net), .MSSIO21_OUT(
        D_MSSIO21_OUT_IOINST_net), .MSSIO21_OE(
        E_MSSIO21_OUT_IOINST_net), .MSSIO20_IN(
        Y_MSSIO20_OUT_IOINST_net), .MSSIO20_OUT(
        D_MSSIO20_OUT_IOINST_net), .MSSIO20_OE(
        E_MSSIO20_OUT_IOINST_net), .MSSIO19_IN(
        Y_MSSIO19_OUT_IOINST_net), .MSSIO19_OUT(
        D_MSSIO19_OUT_IOINST_net), .MSSIO19_OE(
        E_MSSIO19_OUT_IOINST_net), .MSSIO18_IN(
        Y_MSSIO18_OUT_IOINST_net), .MSSIO18_OUT(
        D_MSSIO18_OUT_IOINST_net), .MSSIO18_OE(
        E_MSSIO18_OUT_IOINST_net), .MSSIO17_IN(GND_net), .MSSIO17_OUT(
        D_MSSIO17_OUT_IOINST_net), .MSSIO17_OE(), .MSSIO16_IN(
        Y_MSSIO16_IN_IOINST_net), .MSSIO16_OUT(), .MSSIO16_OE(), 
        .MSSIO15_IN(Y_MSSIO15_IN_IOINST_net), .MSSIO15_OUT(), 
        .MSSIO15_OE(), .MSSIO14_IN(Y_MSSIO14_IN_IOINST_net), 
        .MSSIO14_OUT(), .MSSIO14_OE(), .MSSIO13_IN(GND_net), 
        .MSSIO13_OUT(D_MSSIO13_OUT_IOINST_net), .MSSIO13_OE(), 
        .MSSIO12_IN(GND_net), .MSSIO12_OUT(D_MSSIO12_OUT_IOINST_net), 
        .MSSIO12_OE(), .MSSIO11_IN(Y_MSSIO11_OUT_IOINST_net), 
        .MSSIO11_OUT(D_MSSIO11_OUT_IOINST_net), .MSSIO11_OE(
        E_MSSIO11_OUT_IOINST_net), .MSSIO10_IN(
        Y_MSSIO10_OUT_IOINST_net), .MSSIO10_OUT(
        D_MSSIO10_OUT_IOINST_net), .MSSIO10_OE(
        E_MSSIO10_OUT_IOINST_net), .MSSIO9_IN(Y_MSSIO9_OUT_IOINST_net), 
        .MSSIO9_OUT(D_MSSIO9_OUT_IOINST_net), .MSSIO9_OE(
        E_MSSIO9_OUT_IOINST_net), .MSSIO8_IN(Y_MSSIO8_OUT_IOINST_net), 
        .MSSIO8_OUT(D_MSSIO8_OUT_IOINST_net), .MSSIO8_OE(
        E_MSSIO8_OUT_IOINST_net), .MSSIO7_IN(GND_net), .MSSIO7_OUT(
        D_MSSIO7_OUT_IOINST_net), .MSSIO7_OE(), .MSSIO6_IN(
        Y_MSSIO6_IN_IOINST_net), .MSSIO6_OUT(), .MSSIO6_OE(), 
        .MSSIO5_IN(Y_MSSIO5_OUT_IOINST_net), .MSSIO5_OUT(
        D_MSSIO5_OUT_IOINST_net), .MSSIO5_OE(E_MSSIO5_OUT_IOINST_net), 
        .MSSIO4_IN(Y_MSSIO4_OUT_IOINST_net), .MSSIO4_OUT(
        D_MSSIO4_OUT_IOINST_net), .MSSIO4_OE(E_MSSIO4_OUT_IOINST_net), 
        .MSSIO3_IN(Y_MSSIO3_OUT_IOINST_net), .MSSIO3_OUT(
        D_MSSIO3_OUT_IOINST_net), .MSSIO3_OE(E_MSSIO3_OUT_IOINST_net), 
        .MSSIO2_IN(Y_MSSIO2_OUT_IOINST_net), .MSSIO2_OUT(
        D_MSSIO2_OUT_IOINST_net), .MSSIO2_OE(E_MSSIO2_OUT_IOINST_net), 
        .MSSIO1_IN(Y_MSSIO1_OUT_IOINST_net), .MSSIO1_OUT(
        D_MSSIO1_OUT_IOINST_net), .MSSIO1_OE(E_MSSIO1_OUT_IOINST_net), 
        .MSSIO0_IN(GND_net), .MSSIO0_OUT(D_MSSIO0_OUT_IOINST_net), 
        .MSSIO0_OE(), .REFCLK(Y_REFCLK_IOINST_net), .SGMII_RX1(
        Y_SGMII_RX1_IOINST_net), .SGMII_RX0(Y_SGMII_RX0_IOINST_net), 
        .SGMII_TX1(D_SGMII_TX1_IOINST_net), .SGMII_TX0(
        D_SGMII_TX0_IOINST_net), .DDR_DQS4_IN(GND_net), .DDR_DQS4_OUT()
        , .DDR_DQS4_OE(), .DDR_DQS3_IN(GND_net), .DDR_DQS3_OUT(), 
        .DDR_DQS3_OE(), .DDR_DQS2_IN(GND_net), .DDR_DQS2_OUT(), 
        .DDR_DQS2_OE(), .DDR_DQS1_IN(Y_DDR_DQS1_OUT_IOINST_net), 
        .DDR_DQS1_OUT(D_DDR_DQS1_OUT_IOINST_net), .DDR_DQS1_OE(
        E_DDR_DQS1_OUT_IOINST_net), .DDR_DQS0_IN(
        Y_DDR_DQS0_OUT_IOINST_net), .DDR_DQS0_OUT(
        D_DDR_DQS0_OUT_IOINST_net), .DDR_DQS0_OE(
        E_DDR_DQS0_OUT_IOINST_net), .DDR_CK1(), .DDR_CK0(
        D_DDR_CK0_IOINST_net), .DDR3_WE_N(), .DDR_PARITY(), 
        .DDR_RAM_RST_N(D_DDR_RAM_RST_N_IOINST_net), .DDR_ALERT_N(
        GND_net), .DDR_ACT_N(), .DDR_A16(), .DDR_A15(), .DDR_A14(), 
        .DDR_A13(), .DDR_A12(), .DDR_A11(), .DDR_A10(), .DDR_A9(), 
        .DDR_A8(), .DDR_A7(), .DDR_A6(), .DDR_A5(D_DDR_A5_IOINST_net), 
        .DDR_A4(D_DDR_A4_IOINST_net), .DDR_A3(D_DDR_A3_IOINST_net), 
        .DDR_A2(D_DDR_A2_IOINST_net), .DDR_A1(D_DDR_A1_IOINST_net), 
        .DDR_A0(D_DDR_A0_IOINST_net), .DDR_BA1(), .DDR_BA0(), .DDR_BG1(
        ), .DDR_BG0(), .DDR_CKE1(), .DDR_CKE0(D_DDR_CKE0_IOINST_net), 
        .DDR_CS1(), .DDR_CS0(D_DDR_CS0_IOINST_net), .DDR_ODT1(), 
        .DDR_ODT0(D_DDR_ODT0_IOINST_net), .DDR_DQ35_IN(GND_net), 
        .DDR_DQ35_OUT(), .DDR_DQ35_OE(), .DDR_DQ34_IN(GND_net), 
        .DDR_DQ34_OUT(), .DDR_DQ34_OE(), .DDR_DQ33_IN(GND_net), 
        .DDR_DQ33_OUT(), .DDR_DQ33_OE(), .DDR_DQ32_IN(GND_net), 
        .DDR_DQ32_OUT(), .DDR_DQ32_OE(), .DDR_DQ31_IN(GND_net), 
        .DDR_DQ31_OUT(), .DDR_DQ31_OE(), .DDR_DQ30_IN(GND_net), 
        .DDR_DQ30_OUT(), .DDR_DQ30_OE(), .DDR_DQ29_IN(GND_net), 
        .DDR_DQ29_OUT(), .DDR_DQ29_OE(), .DDR_DQ28_IN(GND_net), 
        .DDR_DQ28_OUT(), .DDR_DQ28_OE(), .DDR_DQ27_IN(GND_net), 
        .DDR_DQ27_OUT(), .DDR_DQ27_OE(), .DDR_DQ26_IN(GND_net), 
        .DDR_DQ26_OUT(), .DDR_DQ26_OE(), .DDR_DQ25_IN(GND_net), 
        .DDR_DQ25_OUT(), .DDR_DQ25_OE(), .DDR_DQ24_IN(GND_net), 
        .DDR_DQ24_OUT(), .DDR_DQ24_OE(), .DDR_DQ23_IN(GND_net), 
        .DDR_DQ23_OUT(), .DDR_DQ23_OE(), .DDR_DQ22_IN(GND_net), 
        .DDR_DQ22_OUT(), .DDR_DQ22_OE(), .DDR_DQ21_IN(GND_net), 
        .DDR_DQ21_OUT(), .DDR_DQ21_OE(), .DDR_DQ20_IN(GND_net), 
        .DDR_DQ20_OUT(), .DDR_DQ20_OE(), .DDR_DQ19_IN(GND_net), 
        .DDR_DQ19_OUT(), .DDR_DQ19_OE(), .DDR_DQ18_IN(GND_net), 
        .DDR_DQ18_OUT(), .DDR_DQ18_OE(), .DDR_DQ17_IN(GND_net), 
        .DDR_DQ17_OUT(), .DDR_DQ17_OE(), .DDR_DQ16_IN(GND_net), 
        .DDR_DQ16_OUT(), .DDR_DQ16_OE(), .DDR_DQ15_IN(
        Y_DDR_DQ15_OUT_IOINST_net), .DDR_DQ15_OUT(
        D_DDR_DQ15_OUT_IOINST_net), .DDR_DQ15_OE(
        E_DDR_DQ15_OUT_IOINST_net), .DDR_DQ14_IN(
        Y_DDR_DQ14_OUT_IOINST_net), .DDR_DQ14_OUT(
        D_DDR_DQ14_OUT_IOINST_net), .DDR_DQ14_OE(
        E_DDR_DQ14_OUT_IOINST_net), .DDR_DQ13_IN(
        Y_DDR_DQ13_OUT_IOINST_net), .DDR_DQ13_OUT(
        D_DDR_DQ13_OUT_IOINST_net), .DDR_DQ13_OE(
        E_DDR_DQ13_OUT_IOINST_net), .DDR_DQ12_IN(
        Y_DDR_DQ12_OUT_IOINST_net), .DDR_DQ12_OUT(
        D_DDR_DQ12_OUT_IOINST_net), .DDR_DQ12_OE(
        E_DDR_DQ12_OUT_IOINST_net), .DDR_DQ11_IN(
        Y_DDR_DQ11_OUT_IOINST_net), .DDR_DQ11_OUT(
        D_DDR_DQ11_OUT_IOINST_net), .DDR_DQ11_OE(
        E_DDR_DQ11_OUT_IOINST_net), .DDR_DQ10_IN(
        Y_DDR_DQ10_OUT_IOINST_net), .DDR_DQ10_OUT(
        D_DDR_DQ10_OUT_IOINST_net), .DDR_DQ10_OE(
        E_DDR_DQ10_OUT_IOINST_net), .DDR_DQ9_IN(
        Y_DDR_DQ9_OUT_IOINST_net), .DDR_DQ9_OUT(
        D_DDR_DQ9_OUT_IOINST_net), .DDR_DQ9_OE(
        E_DDR_DQ9_OUT_IOINST_net), .DDR_DQ8_IN(
        Y_DDR_DQ8_OUT_IOINST_net), .DDR_DQ8_OUT(
        D_DDR_DQ8_OUT_IOINST_net), .DDR_DQ8_OE(
        E_DDR_DQ8_OUT_IOINST_net), .DDR_DQ7_IN(
        Y_DDR_DQ7_OUT_IOINST_net), .DDR_DQ7_OUT(
        D_DDR_DQ7_OUT_IOINST_net), .DDR_DQ7_OE(
        E_DDR_DQ7_OUT_IOINST_net), .DDR_DQ6_IN(
        Y_DDR_DQ6_OUT_IOINST_net), .DDR_DQ6_OUT(
        D_DDR_DQ6_OUT_IOINST_net), .DDR_DQ6_OE(
        E_DDR_DQ6_OUT_IOINST_net), .DDR_DQ5_IN(
        Y_DDR_DQ5_OUT_IOINST_net), .DDR_DQ5_OUT(
        D_DDR_DQ5_OUT_IOINST_net), .DDR_DQ5_OE(
        E_DDR_DQ5_OUT_IOINST_net), .DDR_DQ4_IN(
        Y_DDR_DQ4_OUT_IOINST_net), .DDR_DQ4_OUT(
        D_DDR_DQ4_OUT_IOINST_net), .DDR_DQ4_OE(
        E_DDR_DQ4_OUT_IOINST_net), .DDR_DQ3_IN(
        Y_DDR_DQ3_OUT_IOINST_net), .DDR_DQ3_OUT(
        D_DDR_DQ3_OUT_IOINST_net), .DDR_DQ3_OE(
        E_DDR_DQ3_OUT_IOINST_net), .DDR_DQ2_IN(
        Y_DDR_DQ2_OUT_IOINST_net), .DDR_DQ2_OUT(
        D_DDR_DQ2_OUT_IOINST_net), .DDR_DQ2_OE(
        E_DDR_DQ2_OUT_IOINST_net), .DDR_DQ1_IN(
        Y_DDR_DQ1_OUT_IOINST_net), .DDR_DQ1_OUT(
        D_DDR_DQ1_OUT_IOINST_net), .DDR_DQ1_OE(
        E_DDR_DQ1_OUT_IOINST_net), .DDR_DQ0_IN(
        Y_DDR_DQ0_OUT_IOINST_net), .DDR_DQ0_OUT(
        D_DDR_DQ0_OUT_IOINST_net), .DDR_DQ0_OE(
        E_DDR_DQ0_OUT_IOINST_net), .DDR_DM0_IN(FIC_3_APB_M_PADDR[30]), 
        .DDR_DM0_OUT(D_DDR_DM0_OUT_IOINST_net), .DDR_DM0_OE(), 
        .DDR_DM1_IN(FIC_3_APB_M_PADDR[30]), .DDR_DM1_OUT(
        D_DDR_DM1_OUT_IOINST_net), .DDR_DM1_OE(), .DDR_DM2_IN(
        FIC_3_APB_M_PADDR[30]), .DDR_DM2_OUT(), .DDR_DM2_OE(), 
        .DDR_DM3_IN(FIC_3_APB_M_PADDR[30]), .DDR_DM3_OUT(), 
        .DDR_DM3_OE(), .DDR_DM4_IN(FIC_3_APB_M_PADDR[30]), 
        .DDR_DM4_OUT(), .DDR_DM4_OE(), .REFCLK_0_PLL_NW(
        FIC_3_APB_M_PADDR[30]), .REFCLK_1_PLL_NW(FIC_3_APB_M_PADDR[30])
        );
    BIBUF DDR_DQ8_OUT_IOINST (.D(D_DDR_DQ8_OUT_IOINST_net), .E(
        E_DDR_DQ8_OUT_IOINST_net), .Y(Y_DDR_DQ8_OUT_IOINST_net), .PAD(
        DQ[8]));
    BIBUF MSSIO3_OUT_IOINST (.D(D_MSSIO3_OUT_IOINST_net), .E(
        E_MSSIO3_OUT_IOINST_net), .Y(Y_MSSIO3_OUT_IOINST_net), .PAD(
        EMMC_DATA1_SD_DATA1));
    BIBUF MSSIO26_OUT_IOINST (.D(D_MSSIO26_OUT_IOINST_net), .E(
        E_MSSIO26_OUT_IOINST_net), .Y(Y_MSSIO26_OUT_IOINST_net), .PAD(
        I2C_1_SCL));
    BIBUF DDR_DQ0_OUT_IOINST (.D(D_DDR_DQ0_OUT_IOINST_net), .E(
        E_DDR_DQ0_OUT_IOINST_net), .Y(Y_DDR_DQ0_OUT_IOINST_net), .PAD(
        DQ[0]));
    OUTBUF MSSIO17_OUT_IOINST (.D(D_MSSIO17_OUT_IOINST_net), .PAD(
        USB_STP));
    BIBUF DDR_DQ6_OUT_IOINST (.D(D_DDR_DQ6_OUT_IOINST_net), .E(
        E_DDR_DQ6_OUT_IOINST_net), .Y(Y_DDR_DQ6_OUT_IOINST_net), .PAD(
        DQ[6]));
    BIBUF DDR_DQ1_OUT_IOINST (.D(D_DDR_DQ1_OUT_IOINST_net), .E(
        E_DDR_DQ1_OUT_IOINST_net), .Y(Y_DDR_DQ1_OUT_IOINST_net), .PAD(
        DQ[1]));
    BIBUF MSSIO11_OUT_IOINST (.D(D_MSSIO11_OUT_IOINST_net), .E(
        E_MSSIO11_OUT_IOINST_net), .Y(Y_MSSIO11_OUT_IOINST_net), .PAD(
        EMMC_DATA7_SD_VOLT_CMD_DIR));
    OUTBUF MSSIO34_OUT_IOINST (.D(D_MSSIO34_OUT_IOINST_net), .PAD(
        CAN_1_TXBUS));
    BIBUF MSSIO25_OUT_IOINST (.D(D_MSSIO25_OUT_IOINST_net), .E(
        E_MSSIO25_OUT_IOINST_net), .Y(Y_MSSIO25_OUT_IOINST_net), .PAD(
        USB_DATA7));
    BIBUF DDR_DQ12_OUT_IOINST (.D(D_DDR_DQ12_OUT_IOINST_net), .E(
        E_DDR_DQ12_OUT_IOINST_net), .Y(Y_DDR_DQ12_OUT_IOINST_net), 
        .PAD(DQ[12]));
    OUTBUF MSSIO31_OUT_IOINST (.D(D_MSSIO31_OUT_IOINST_net), .PAD(
        QSPI_SS0));
    
endmodule
